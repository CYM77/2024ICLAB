
// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
M-CX5[;(TP#W^@U/J#R4LC@/W0O7GgZ<57D,DG3XD=J>.PT-f^6d-)_49(X]=335
5F,beD2PP@MIUed=1fXTZOZ&a&[G#8fO+N<W+^U5a<9V5,)1@H;]OIeH?eEZaB\b
/d=UD#a_;@?U\H@G9Y_/(>X\?bD1;/g&^5]bII&]NFHdZL;_J>[5eR.29]#:2IZ_
U?DROU;A2<=2+H(Y:gQO0M4G\.[Z4=J>DK8X9g[J-]C1^eH+Z4Z&Q5>&A42O4:cL
/#880;G=+4B/)L/3AcA18-L>P\3cZ&&D+\J#W9<YDdH&^EI&b)M/+?Ge2#@8>S]Q
-aAH3](Q-JUD8b<dTe7P1JS/e?1KeBbK++aGCYS#,>c\#2EG)?fWeCVN15H<A@I:
43,_RePD-A,Te]2?A0Za\U?&W@a<8KaK+4.PB5WVZPEYEOV4(>()/;b.KK1Lf>S3
GIF6ACYF,#gAYC2H\K=VKA&f>)Y,MIK^3KT90gV++De7(cdd&]R?@<b&S)a(c(9L
S<X:SZ3F+Va<G7&;)ZT=3&)gET1,fGS84>OQ2fA+e8aGYI0NZATU/AE<+?N)e10&
L#Z0g7[4>>K/AbC99dXJHU#)PMPH^3Ta?LD>ZPeIFWLQ^)0A481)P+fHDOQ@&g+/
,),+LQ;L0D<]#>SDHP5NXKHIL?+1B71eBeH3RXAN.WC9EITCV\8V[DB/UI@XQBX)
?]Y[#8@7Pe6/3.e+EfPMR-Z8dY5<W<OP\9AQ7?;XgfK\>bb+P2VTGEAM6WNB:E4S
><-/U7K>2LZJZ1Jb8b=Z,1A:J&.b/TAJ:1(I;c;?,<^_<EcQ0#MQH5#f/#AY7gaO
]dc-J:6J]a1:6IfE^K=M>bJ(08XbIJa,-4gSPANEB.E_;d#YU[=O[(6Z9^TM>QYX
Td,7E6QVY66HbK//:=-4BD7MEN=fYF[&5F/G.RY7E(@=eXP0[6L1;4.93E:?Mf6b
,D<gDI::CeP,0b&L4b^?e=IA<_260XGRK26;??#D)A1M;?Mgf?\>+A2K.7KZUXT=
L=WN6X\,<(bTEJ9.[].Hd(G_\FPeFS+QZ-9RXeg2YL+C<W0:-2#5H31HfR?[?+]N
)0PY)PfFJ8g_=FJE<N2Q7KN:aELQ5:_BVSeB39X_4D-C_>1d9,?HUF_W)8[)S16I
Y50]7Yf,]=(324]<<S=#Sf6bDbR]U^g]#9ZP=C^3H:W7gUNfW<bOTBX19-97ac\(
SG[T-gB:TZ20)TdPO8@+bfgZ;>b9Wf]agL;I4:#<T<KY[5R9]DM#Z>;5T[c@:(aS
JX(YRXA:2+)TR24DW3N#7IfY>#H1D]L\XMEVEUF8)eX4]WSI2N<HW^=OB^,6,BH4
_ZQCUcb]D?0NJ)C8a.#)HTKG8LGX3NMa#1_g+WIdJ74Q(3Fg&5?6L4Ig\fR.[AS2
#RT;W[29X+ad<;e8TCIN[.9g<CZUJ&?_BRX[99P=\??c@DCf4J9U1T&VCCL?Pf2M
><>Ab6fJ,b]WbO8Q:g\3d?8=EZLbFdRNf<6<,e,K[CR4G6RPBf/36XPZM_QYGbU1
C3(/D[[GE8f@YMNafYKS1_/T19HR)1-):W6Tb;M^dG_a:AeId0Z(KK9]UL#BR)^M
^H&R9dCRLF-L2/\,La]bE&\MQ8+]X89T^H]]:U_d:W&BQCW<>6)cM]T-\Q+3<]\X
S?/OUPA<.96_]N0&:Bc_Y)\(N[1EOQaQ3<,XEP3XaTf<26J=<N]A>SMN4<N([44Q
/RI&/02=R]J8UV1]9gA19K;9LXV,F)RVEX\,_J?]P@\78>M[MFNDGX69dJ2#B+/(
.?:9:c<>Y=&<;:I]GR_GWWZY.],I08bI2FBDX<6LC_)WP?TYA/M[>FS2U=F9MS]a
11fb)#)^+eW-CHH[Y070>=Q,b<D]UYZ8YJ+b0+g^1acLO(>H]9G];(M0_R9f)gQ]
L)1ea8afEH=<L5\7BZXf?[>Ybed,X>\XabC[8UR&71UE33;#/>5I)/+4C3[bBC@\
Q>M,_gBRTPXTWOVRcXU6XV4NHJ.OQN7c[KNb9:?^c33E(PJBTAIN(DI7D=./3d3X
A\6C/;\cMDP:>ZKI--4DSF(/3-:(J1GUMP:VJ^.Tc8T0L+>cX^PLV?@0O0BL=YUJ
+g2I#[f2V^+F4UYa1@7QXM,NcQ.XEF1gOdEOMFO)Efc19-gdFG_@0D:]EdN(DC5#
L]\?K]EQJA^\\5_5#fe)D2-c^ESOPGY(W_\KJQI5MH8P_DMc>f//6e_c@;V-E<df
ea7-;A_dGM0a\:)CI+IbgHJH6RM:f?g[;1,:aOS.SZT18I3fLg&DO61@;(G6>J\L
W4UG@\(>I.Be-2DV(?ge^D@^M_&JE)g^-7Qd^(;_5UKIJ//LK38+D3RO\\.IATHW
L7=[/8LgRIR1^R71:>>;)@7;\=?+()O1GPFMK)1N-8U5,;@^Cb^0C#3AYL]9YS=:
Z>4U7JF^D8G^3O#;9Ua^,5?Z]PK_gT\34bBN\I63/;D.XEdR9Q2D1RJI;La\,T?)
)9KM0>A8QI)UHC,R3YK8G#GK^<SgL.&IVTcIQM:R&af>1FKO+HG=a=:8:4:b[^H3
G5=2;RN2HB-/C)/de-LJY?f,&,_5b6_8[SAZ\8P;L9f3?_=B:?&[/Z2F7Td.ZU/D
GXb1DdEdXRDD/X)C;/IIR/_]Fe=FBX6C,^P0N8fSHd(/XFA(0&_X]\A;PT./2/-5
<:F_IbFUQ<_R=S+\Z@TU>:dZ,R5P4#)/AgTEI/dbB6[:bKC#:-O4>C^#e/#F,:F,
P/O/adIH<2T]OZe(EFWNY24@KQLeJP=<XEQA?5=>4F#+5SNEgZWDTQS12JIY>]\N
^K<eO@@QN@dPU]K(AET2?NUKH7g1@-:.Z-d,J#YP3>HN4:F#[+6DH(H=>?,Z0Kde
<#5KHgPP?>X3YWM-L_PcKGZ?)1Z3I1[P1c#K:NfIW+EP</UBZEEQ0^e],3HOS4XX
R6cST8E/[_.\1>g&>7U3SL>1XET)c8Y.^1N]W+>TJS=-^AQG3N(A#4)RP#>(Zd-c
.d1F[^4.7SNae=)C42WD0AP1HLEf]EVXO/8,H=T[V?-Q1GYQJ#>e61QKSB=]ZYCT
M#>FU:Ag#W1=3L@eV:Z8ZJ71dTNfA3N5cM9ffc7JB&-2VLMZZQ]=(JY30<5;>c6V
Z5S/<D0M;e:g3>L;g[cH46IDZ5W?G]85HZR_BIccRf);gC_JO5+MW=,=c.+OYKaG
UeH5Rge7(-c]RBNZR(R,2Q(_9(_Q3N3,[cS;4HB&E5L/QA06\[9.9TEMb1Y=S[5B
;-X546K;a[1,?(:AA3?PTB]@D9LH9&6SQ#ca<:2,M+YI0TdOMObU[+]ZZ+>56.d(
;Q\M<VKS/gI,DQ6.I.aTaJ(#4?e2W=KT<ATLgLXR<2O=?V5WI4F+3)-V0;_]U&H+
=CZ;33Y?S:J:P4KUf.fc233GE<ZQK^\a\)<8\I(S]^=9eWe<Y>eVXE3)TcGS:?D_
&)EaJ;eMJZ7WE7YcHW)0,\RAXfW:ScF3E#-K],+B5.:=@>EcH1E]<&<d1BcJDV5W
[Ye&CL28&M.@QWCN<^PTEeV9F1)fIC,Ng/c]&Y5FGG.D^S+.7BI(0AY;+42(]Q7T
-[(RUg&-WS5R0YV(8A1b_S.WP\Y-bDLA]JTe0=E=(RE@X9-U-;-?g.BK@geJ5)(/
ZWIX5U+-PQd/B1=(XU?FTPP:5bHI2ZP1cR+d5R?<VV1cS\JS?=/4&H=?W:e@DfFG
VfLD8@E0&^G2:U&aD7UXeM;)LW&KL&09&1IBMHQ+:)[/W?EVX_+TF;Z&8ZB&0\1W
@e,5c6JOX@9XAW()43aIEJANWGF+FPPe7e?\7W6U1^.SVdGH07Qd#cI:(?2S<H@D
cW1X9L^K?DS9#:V28d,J.M]^]M;GH\7<TSPcDRHO58fQ+6\4;/e22+NBce0F=B;H
<HG&NAH+#P-5e@^eS]Y8;5ZC91[41_a/-=EIWeV;R=VIaSG0<g.601RRK_HWU,e#
Sc5L56KF66P]7a^449RS3.WPMXLD>=-9OP=,01//3&1[-A>KX03NQfYO:aFO^ON-
=GA2GSQZ?^U7W&Vb#0<&F(:-LMPW?CDRN_6D59Ag>EU.M9e4<)@Y(+]L71QLa&#E
D.dcGf(F=2OAGVDc+B[I/K1/4+3Lg4K<:0ICX.\HT22YD<aa13HI@+]HZS._)3ZO
ac#11Q+/#5:9Qd@0+d]32#c0BWR(.HDA6\\?AW)<(Q&69R@?#K7ILL;aT1Sc6>c>
P=O&EN,+ad<TeS86#F;B(R+/#@cg/?X@4cbRcG#a@AW<U_07cVAS2;VbII]-f5I=
A,NMMW:OP/0<\gg0A29=AfO7:M?R5]5=BCa&GH3BN/I0>N7dYfWW>C[^X-;C?5=P
[4e7(.=VVN5U0\BST4=]E+R>#8a,-GZAbAO,TAY^(ESf^:9PQMI84Va3TN68b.:c
[-TE0V66#.=?4,[E6F/(]Hb7=:Hb6_<PF2E\)dF4[?U,MLVL,DYEJ[dEEK0_dRfS
7@=_E-VZHgfSKg4W0(aB4g_Qg#<c5I45Z-B@MGF4Wb_CbF4(#Ad)e0T73VAfO)XJ
/4?;ZTbWPF0?8N-&P@90EP,?=;d.\NA0ZM9AL<a_<:Hg.35_4BBO^R&DbEW;4(35
;Q,JD9FB<T2I5e-E]&,-[f&WYb1<#16>;[43OJc8:g?Jg1>(D(SWNSK-[OJK25M+
L,cLB>:&eV7Y>K,][,)YFLHDU3X6)IMDd=S97N_5,Y.>)?RQM?[A:@c-J0+eU>Va
F8UgNIYF.Y+;Y-LR5-e;eIG60.41W4FDADIZ/JBf4e-<dIB?g1M<TU1K(E0]]9@P
QKaV#TLRL#GARHO,;B8YV4=P<1,CV=E9DNM-CG4:EWCe7+OCQ^.&]0HLUNPKg7/P
A:[-LH)Ub]H4HSg5XZ<GIAP)@7J3dggV.9a)0V>P>^3JJASaDC0a;,dY46G<Qd)J
<D@S(/ZgTE24O#7I&6fUN.1TPL@WB1AJ4WBCMM6)c]HL@E)D0@8c[K[<4U#:NGZV
8C+I^;d_4RQZ@c62-=[]KHY.dX^6(UC1g&I@#1F-^>KZ/gIR]E9-2@JSRd\?<?G-
E(;5[F@NSD;SY?:WHd#,gCGBaSJZ9C\Vf\V/@9UZOM-=g<&SSZ@B)9.E+14FA,U#
AIDNeJK-RbS+UCUWX[_Lf[HIET@(9S1eFU[W<SJ1fA(VG<MNZ1M^XXM6&WD[YTFG
)a\2bWQT-SE=\1NO+QBJC_Xg;eZAKfe^.PI@TD&G-gU18Z\E>AK7P,\VBSfBU+@1
?E.2]7Z=;NN?^BHR?M[TEIOBEG\JeS85?X>d1OCMGc@0PM7F46OF+;-aG[2R^[IF
6)LeB.=[>MG\&E54@_CA/FHaLbQL#FGaF7^^U1^:b7]g,X5G@9?g^)&46@YBL.bO
eLG@ZXK;?-2VAZA&beQDVAg,WB#XReEGU7SY6ZP7;^L\.Y>;X2)fO6AKQLB9)LK[
&H3W-GgMRF[7&L98;4dVc)5B^E8B]GCR3\.WU?)F1C[e/99G0CA:?/[c>;O6HLeN
LfW^a)6EL?cAV4Z=GJW]D3@GUZN][,.TecBX,[a3TYW+]XD\8LYZI_3c,26T0f]1
(VG\,SRS48_N/-MWdJB7&YLLTe0d[7cX+\M3,\C#-]P6,Y6,AN&V^IF0K6GUf6H1
@e]9Ke@BJ/\EIf+F-V62]1BGbC2X3RY>WE27\^[WM9,I9fL;c/;FA7Oa.4,<FaAJ
cRR1W>>1eMB:V?R0L,dg(IdM41AcM6.:P^NcR=/I1.?25)cfX5@H7[X#:/HHf^#)
DEL6^KcM[OVY\+12,G(e@<abf#OQ<;FLS@+K:7&T2T?Wf-:==LY_01P+9P\0aQNF
X5a5fB3YVBPQY-dTO3dLJN+GVIc?U/AUW6[W6+YVY80=Z8>?cYT8U8]I4F]9L5Q&
)[66JQ],D=2]<155VdS>#.e,FOabS@0KSJ6,5L]>.&?YTd.QD03>7cFP3;/J7ecQ
1dMeT]^X&H_U.g-ZJYT/7<6f:#bSA^G@+aG/-,>L(WHAM.,B9fT//<J?gMO9G+e6
S\O9YA^>7a1QN?K.@S(a25@APYD)f;_9)6<&3H-Rc2C9(Z>/FHZ>>c_><=610eOJ
P>]U<dGTD3RKfG:fNd(K\dYaK\=_)>g]5(.MO1C2/(a&\+L0B#5(L.VCUQQcfTQe
fLIYI1PJX#+X)V9:c?C_,3KR<DKf5-HW:/9DUCM^0LDO9PL+?U+P?FNGaV_);\>L
7acHW?0;Y):V7A9I3f[Ufe,P5C1#c,^J.IPf/,+91NZa0\&NccBHI5,3H+b7C)HD
:GS3C?.#F1Of?fLcOQ>[BAJ43F4OQTTa&&58e.:4UB\+/H0&7fYGK_dLNA?7Y</a
-f)>+39MZ&E?+,gB9L@;:ASU3aE5X#L]J;AOe@5J4LcT&I<E]<+IBWfeTd8O#4VC
SdUOGR-I(73<b5COKZ,V[8,;f],=S8J@I1addQ,9;R(7Bd&2[TL0:Y[:c3I]-N6C
.OPCKK6SL,[##2EgZ=1JW8,fbT<7bfKPL+@HA,7Y5]\,cPVU&6<#UKJ=f2c(3X>.
YW3L?FAO_B@>:3aP=>)]((<XM^2b++[YS6M]6#HDTT2#4\=+QDe>TB=aa6XLf[dK
DT/=B.bDIV\Qg5?7VF:F#V.QP78Y7SP2@e>Ef58@]JaD\;EY=ZK4X&e<95]A.CQC
(^fRIU4AL+34f>d_J(9^@?L6NecaRSXc43aHdI3MU^Af64MCdXY8E-GDg#\CEW</
Y<XRX+7Xf\gO=(C35He&F6g/Xb[\]:DBYDG:+_+b(aR0:91bBS45Nf^,SZ8N6@/b
KB93.XS@FJ8a;E:e^Rd^6=O1N#WJg/=BGZ??d:Pb7=Y(fgcEH.AdNZQM-+(N;6U_
GU5@[,CMec:L.e]Rc@;+ZEXQ4:)_,fJaA#eRL/)UD=I=S2B5-B9DLeX>W\e4Z+Z7
[\TA_<T@ZX0,N()FFfWKIcWOSeGQU,<3f/7#39c^(L(O/N5?#3ZBN.0A//d6Z+PY
EFWW@e,)(]5^d(O^1TZ4fO&8.BQMJ9;3=33()D>(2DM3R3ba7Wg\B:5B+7MHR9^5
8,)ID?=]INc=4;V^=<YJ+QY(B,=IFA&aFFf2,;Z.(#5d/O3;U;Jg9D)3=a.5^>af
DR]5cg-1I9NNe1/3cWD/)E<b-Jc34GHO\>A#.O5C^#3+&\D==Q9EF_>?([7]3TVH
Yfb/B0e)A/HD:&AMbES9Hf\]S2b>P\dP/B=:Pd)K>4,3Z4JR5[1e6\4-T+/_6123
8]FJQK\ZVN<@+@^MU0c:E<LKg#c;1XS39.WO=KP1/J<&eZG[MJ:2MT0Pf(OX]9I4
[e#BCN=Hbc(\P\.>B[E[I,ICI?QV0\GYF6_dW[M1cM3=BZg<WO#Z2O#E#J2@7L5=
F#L=/=]0g6>aK[\LFL3G+;TgUM6-;0),J@Z+MK[,K+O\dI:8M\e,YKLf:cTc;9\W
fFbbdegX=:GaM4W@>7R>\8)@2cTC:WKD._F=)@0AJM,:?M.(G#7)7<L^5H6QZVA&
CfbLgdg3L/Sf\@IR)5X.+4)@WA)E6VSB@89QW^37>:MEU)PB/.Y4,G[[4bcaG::6
-:Y\\e6Q-1\NYN;TG\NC4BdbKY4G<a@T<6F41^UTfHF7JL;OQYA)U1<RM&EIG+ga
VWX2_I8MRMI05NUFJVSK7NSV5G;P14Q9TPAJe#11W/2GV/(S/NUXIP3OV#PZ0?VW
8\7a-K1-[/S[6=<R\078Of([=a-5<Kg#JJZG2ZdM)_b+Jb50\F:T_&Y:d<3FA[-e
X4JY+>EV:9&<PPc_ZKZgIEI/>5QX3_FeNCJ]L+N3aF]UD7cCX8)=TOZaAdKOQGMa
7B:@L:(FM/=BXE6@X+Yd.+aJCF8>WO&=XdF25O[g_7Od0<d_88)9eHa^BGE+PCIF
8RVLA\HY3KKX_d&L5RX/=DFI#/-DOf)R27UVK61;cXZV#KTZP;]eF5P\NI^baHSH
@HYa&?_e_#F0E_=XVZ2a<4X87&52b_/,QN_VYQBA/B(Wf05O&G,,&.Ye]@;cD2:>
,.V(0g_8=-L(U),<d)T=XdZe:@2G((L,5<fQ1+H-]AT)=D]0<gO_?9eWM3^G(@&>
?0a?>OE=SE:Qd3J_LA>.)3^Z3dPgOJJS/XK\6:+T,2Z-TK4R@1WJTZ-0+e4GGWAV
+\01;#1T>^2)Tb_++;V^[HD+)0X)O]]L>.9d]I1-0fP0B76H3(0??ZBbWN<5RcLT
L/[N56DaHJ]V]Y@c_3OS;C8ZGNB3AP4Bc08VET&688L^>[+@d?/AD_#Z<7DB1M@2
C-GOJM6?5IFV)Sa5=B0d6M6Tg9?#+E:P_MS:fT2=)T5)F<;c+9\;a>,)#gRB3>A@
/JVB8))F\G=HFNC4aZ8DDHUYJ928=T7LDD(Q\4C+KK/<ELf(gS;(I]/SI6N4Z>cF
?\KOCEMUD>-[G;O5eC48Ma+/O0IS89V<f9T/_4GS((OD+T<W8-bF1TD=:>49R;8>
PUUQWfRM(f99@O]ZF__aN2<-f6[TDff:TCQ1R#)>THT;MD]M97V=fL/C-ULYHU2S
82,eH73S>]M&f/RGE):1IRE<4_,D@gB6+))1L(V=L#BM/EL&DH;Q8@U/IaaKb8G^
[_L/SK9M:)Ua:B:2e:0CD0Z]<R,0_8I8N88H=/CVdYQ4[SL]:b:K?H/VT@M@B\UW
]9de1CVbNf9,(aB07P(X_f+<c&XW:eC<7Q,7.eQLa0#)+OG_<Y-TEfSMU;.U3[5J
V6.C)V70+)&KAg_W@#8c--]3H(2B2SY.LD[c>V#,:Mg-9WBg2_+c_#0YTE6Ta&N@
M@Yc;)E<Ie?O<,WfF-OWQOY<+c)J3CaW=XDEc\W7;L9;D>/UgRBOLAfeML4N-3fZ
+a+CJ+,Y>=3@Q8JBO=29eXQXNNLGJ.G,E[DE,XHDWSIFQf#<Z@DD,aK\g3.;49#H
06)f<eL&O5:A[gR+=VGbIW]5EO\]_F,O0d@73SNd9@V6-VC(<1@(9/DZdEXULgdB
McE=Y]5TcJIUcVK(]0D4Y\30+e.[&:d\dKFOLaDfY8<_e77b5?>d16.J2G#)GY=P
N[O]50^E7^\\L78KOb6V,=c&R=1DgZJV@3EBaQ\.&(/[O+][6HTYHb:60RDP1VEf
fWMSGVK^<0dFG21VAXb60I-b2609A]G6dN\]M.,P=E>::VDZCVV5NN[1QM\L5(SQ
g(GM5T?/R5ZOcY-S/PD_HI9.-+@X=NYK-]HPF]=+X:.B)>eF2DI_=ZPULEL09HCf
<9MPV<#R#H_4e<d>D+eG4cBDS2\7+SWD+O+,1KZ.\@5]gLBBKBXKQdW]NF9bVb+#
6-VEQ-XJfb[?JYTGeWYcAS8fV@982XG+61G>N9:NacN&3AM>\8E-0:dUT(?X-OVZ
R@_+]YWECf&JL\bcU15=-GC.cPN.X\,<6WTX.fMON?HB0&+YgF7(BSI10?1fbZg8
>C,L72dYKLH+N-&73^,5OEYX^W@UaK\Y0:a(W)E=W7MNDPC7\WfRI-]E,4?^9N3J
IZ?#=d?^a0]KNS+(\G0gW)C9?JIS.Z-_FLO?I&4<_<R9f;gZ4T?[2DQQGOG?4Hf0
BK_3M[@Z\6C92\(-5@W>R2/69VKTfT5>A>LIYS+W.H_(:#/4:?BZ_Db5F7]L^9f5
bWCM>:-1Y)JbP:2(3W3KL)4?4&)gJ\EU<P4IXE]DHWd[1[,CM:=.6.C1e1MGWR/<
;fN>+N2^>K]=0D2WT13:fV_aB-^G\cWW223MR+[Q6^DC#fK+MY@&V,A;YG<B;Y^2
NE/=H5V6_<>JF[OB#>8gLd-SIG4#CWAc[58F4VF[F^a)7YS<\CR+ZIX_UVTN97^O
[@^7aOGG?9MUPCPW<_]Y6S2N3X8<Bb@=4BG&7;4Y7I=cfbRf.4J6YE/,=X3@=VLL
9fYbAMZba7e^Z)>&#/bYHa=4A_c97F2aQC@J#/>MJ7\0#Ta(OCM^RN.EDBBQ1TdL
?[_Z<8PCQD<&#)4UVC>DO2&gO1HKMU\CDA8R9?F,[<3?OeF?L0&J@NPC@8[:[bb1
.7/?P&9V]IS97&7?A+P\RR_)=+ZMXVcWM7+#?@6707D8Bb<aI1g+J10D5=[<6])(
FVR^7,ND?ZV5c\?3B_W;\+8d99&1#T/6YB_?+=^-/H>L-_E#/EL,,)IA-N2N<-QE
,C5&1Y&3&EP^fR1]D)P++?VL@R::)1>^W8CW?4W:,/O4BR/[c82>BT@TQWE#?NGS
F]0N7Va&XST,Y1.98F>ec)6AFb;+>6^[7Cc#W/a1L.>6e5cR<e^XOLNQ:\eT.a,@
@5^Na<L_^1:4M38NF3L=LN>9YAU#6cH5)-Q>PV7?DQ0(#7#((F\,.A:H#TP_Y[>9
<T:Ec7<ZJfB/LD0FQZ>:W?Udd[)VdFI(JJ=DX\:P2cOOTFA9KEIQ0N]W:,^M-]1g
=;a(9E9a9be^9UWD_aN#ZA8XM_[[PI97cOW7B8^4G6(Y&B.aL8ega@3>0UdWNC_e
#;T5;]B-F)B<,W1Q26I6<,(?2aB[MeUK44bV/@54I9SZNFDPSRCF/CCS/P)>D\D0
bJTNMZ5e.:.M@Q86BK[(6M&?_9,;e=bQ?;9>+Z:Dd<?bU9a&D+HZ86c?UHAg0)9.
[10M]90V(Q1gKP0X5.O]M+AR\?_OUGVG(;(7-0O+>0U;1BENg8F;\6,@cD-W2CVb
(d(6OO1HADA_\/1\Xf3UeI#f-g4IV_2Mc868g([eO?;b6Y6B1ME4<GH1&Gc#PbaJ
#-8gdeI;P8D:G<;VA)8I^#/7E:JY=I@](+T[e)=J#+>f_8FHd(UD1((5J;04P_WQ
BfcV:#;]UK1c#?<UY0M6J8H-4U#90^B_]@,,]b;;)fO^TGRGZe-7X\6<S;:]G?=C
NcE(6bdb#1?G_OQ.@>Hf4(7AA[a3X<:,HaRGO7WYXSNH/IW_D_6McKS<H[H;d?Zb
;5.4_/)N-,>#ESXJ\L[;f9\:C2;g__,)>_RgF8_@Q\^D/UQN0E_1I)8PdR#RFR)e
/&ZK33D0:GX2EE:g/acTK;8/1DAaC@adQ;JUUECdaX]U\Z5_=/M,4JZO)4JFO)P6
GbTYYX81fcB6Jg.?KZcC:WP/8C6(78EfFQ0TRd4_BHf1,8@2<41D0D#\bAF]DWR,
c<N=)Dc_(EP?)1c#K2&COF(c3SLZU<2Be&DZd@;Q4.a>8V_>8_0b]1S&6JW<O-A^
eL/VZ@&JL-15@[8Q7[I6I7a9>)1;c>9=Z?4XY1T#/X>=P<+K0.=)A&.=H\#3gc2B
0R84I-WP77g]b,MASVbT1Zd.>N/95)5:1:Jf_(b-SYI&b<PR)H7Q721U3J[_2>>_
A-O,V&^LXBBV&ZE5OM?42-TEb?@W5fLU.C(CE]C;JZ3T(V,B\84T.+4B-&#F#A^Q
85D]Q,:7aPBZT-bW?\U-D9/2_#MJM4[X?V,f&#ED^WAI?B)H?V\2DD^\fKQ^SBN4
U0A3\F?Oc[2HS_dI_YGC+4.)G0M:9RE,/GU?\7U&+XD2.eg>Z+90D<GJ(E3LG1eS
CdaKR)46g)Afe8cUgZ(b/X^,3Xdc0IMJD^[\ZQ/F+7H^=/BD[HaY\F0:d/CVQCK8
YYNL#:9d#a4AP7?]&RQYJ&^acZNI4?Q(W2GE[LBVN/Mc#X0a1)31@W=X]+c1&@If
;R,#P^&c2TP5JJLMN9DSe_>_26MYa_2IGf;0gc]D35DL5#AgX8Adbeb#/Ta_:c3F
K/9UdKP;cS?57;-;8<I2BZK?X>5J995&#R,XT>RIHRU9ESBH?Q^75]K9VgXdgIcY
W+2KW\CG_8<IP7Z2)bB<Wc>2CZcBX@Z#NIKC0GNbP@<^=;JZ(T.J&.20,[V@0O3V
-K,#BN/?J?5?NZ2&/<T5^gc#V(6@TKPSWQKZ,N[a<X&>9UV<_Yf2fO7b9K=dc3]L
77W0ZWCgMJ#Hb[AQ<[/78bA8/6O4NLD10C#[)f3[I=PB:(OP7A&R+gVD^ML4-HCf
CD+/#,+,?PXD.0QIQI)6BfU[33EZR#DS>H#-.&,8eFI@=?YHO\(d(YRG[UZ>]/DW
T^gf-<[Q2TJcJYW4C+b<Xc.0J=;f=dVc/O@2O-L2PAC>C-0&6DgY4&ecT.S?)cIe
>^3M[We1O6>GNTJ\KPQFV#S#4+V?[=U8e)Y3F4.gM1cA@,?R&W6SO[(T3MTMT\2A
7Z-A33?;(XYZJ-FQF)dCTSJE-B994a2_Ze^D#A;NDD?0Sb56EZDNgP1H7Sa>YVcP
WNeLUg=(dN-:1dK,&9K+?=F:6NcVVUYP#&B#J+K+LY<]fRLITd+fM._#X2Z9MZ&P
D-dV?H[:2VNT-I+]C3NbRST-c6^b5g5A7Q\X,AX&\C?fIUR;8U)b:A#.WBBT6SW1
Pg^ccXeeZ.&P&]gSN;5[4LOcG/71@1I4[]?HN/aT?<UO]9WYY3Y+H=O4)V&Y>JF3
/V^7gVFG(UEaWBe):]EI9B8]))]=:[=RH<KLFPXTWYUfS<bNA)R)eC\9dKUfO9E[
[HE+G8O]bdc)9/T?Xa_<Pd.CND7^(-7O8(X==2L4X^AW+B->-+902b+S,\:6VUfS
VLP@Q]@0^XX-J#Pd9ASMYUZ(@#&W^,(O[J34V)53<cNQ-)-CR3Df(>9?&4bJX@CN
DJB_#H=<4^ST>B[=G&VTLJJAd<:Hb:W0,(/)CRFHcC;EVZ.0/b17MO,2:_cOEJ5Y
3<8VJVXC<Q67c;20c_4V<c^DQX2Z>O<?Ja^eFGKIe/gG\MZC,T#g[/<Q)9UW(d<2
=7T0.,T6_/@Db9/+@Kd:^^_fC=5A_.@&?9(X:O=TW(:M/>d)A_#aZ#>+B7_aHE1T
/4OKQeAX>XS18f6KQ2DB)=#e&LHXBJ9ACcg=1&4),2(UJgT5;Z@<gEA9#2&U_B6>
>Q06=(BAfKe<=>9-.9^Re_;CM9+OMG1)6N0/5)A#gC)(#aNQ&)L#;(JX3;<R?9LG
9#(TSI+.B[PVVf#f98PdIFF_;<E.Je+ZRS@4[d50TMUYUc?@+TV)>BEEP7)8ddHW
8b3_dO:#)7:L6Z5U:YP:;Z973J9,&:H.F;NO;W@?3=3J2SDLES2Nf<<I1M]1DKdf
,YAY+_X[9J^SJ^M>d7P]XGdRJ.gPFbTacQ8ga3S\?@O]+D.4#]H/XLSH9V,B\5a8
<&YHG<bML<d>X9>.BT>e@e0Z#)5A[Ubf4\_)X^eY6KfP8SIGCe>T9ZX&&4;YV5?B
4XGdW&G.M3TeD87N;]/]ZREJ]V[BFYM^YOcBfEf3cT61D_FA-SG;Ug3/S8,T[;B9
13UUX:19dHR]BE+9R#;0dVGPI?L<)//B-?)>/KFFH-MU.W[bDIUU7;a0)(,d=>ge
Q+0N.Y[8fNdP@,G-MQLOWV#1cKU<S,e#[BT3e=2R(5E/?Ea<&U9PJYKIOGSHgC8J
/@5:/HUE5O/_Y8HQRYdNb>C]H/dS\Q5bKa;#2CB/QA8O\\@12(A)>P+Ud)J(<B_0
OEW-F7UJU/;\MRPPHfD\U8e7EF(^A=1+\J>N59.1TEEV.#LE,5eL2<g.AcI)1;Q&
-PZc9^.?L^cRd70:9;Sd)8L<0S6BIdLa3Mc-1?9c^V3fH^,FXPfg1MFPABc/PZEK
JKBI-EbADc1:O^2N4J(S]@g2ZV^gJ)SAKD6\;e&f@_g<g#6T?aU@^8?9f)RWg4&?
KU;@SPa+CaALN,?7Y4AY=RVC_cg9Kc8KI#FF3HO97A7S2VJ6]34._=^AP#D3bTG5
,83H:W5BDIU59daR4N4Q&gIf6E.HGTTcXDR?61]_QZb4W_55CRVA/:+<3AB21Ye-
Y+[&faHD=(V<B]?=HTIT2IUF9SJGZ(<:,@S7AM6HGK6DXWRH<W:0c26]aO,^U9]O
SgM^O3Q=;IVIFf[VJJKWI&X.a96+JB3[g<=NNJ#VegQ6JFIQ9MSU_SR^ePf[?UFB
cKCP()2.+5OA)f7;;+O#gTZ:^/M8=PNZ_N8LZTNd6gFHDM2N]D<a8BNf/(&:a6=<
<JaR^5-EH;#Qa^0O_#]a6dPdD-Db(Mb+bL]U&8-^U<I&E&?f59<\c3ITScJYTM3a
0:[FY47J,\3?ULD90)^eE:d3;4XRYPU5RB9DP5V)4Z6>[\=\Xd0J[R1KeT>,>A/K
fbVR1#6.:>V4;C9_#Qgg^_,deN#J8;0K?fAf=WQXLb##+QH&V,Ib1T^CW_6@C>VJ
130E2254g6?U@Oa^@Xc5O#cgL-1F5,&OVJX_1_6^W&<==\\4O6[-EOad.gg=8DFe
c1\Gc>U4F)^[-V7@_@P?JWBgN>X&Z8U^93INGGQYBgOYJ,RJ.]GMJ/ec&NZNB70P
Uc+<)Z(8^X36MW;=d5f9b=M&LA.6P5U8g>f_W^CNg(1P3.D7D1.@&B:A(TE-[:U<
5&9PQ>4Z/_(b8KM)^CJK5FA2aSLKJ:=_WH_;:^CG]]fD+[<_4YQ06UTBBF[8_OZI
3b_FW7CdZ7Q(D<O4Z([_9Cb:\-9f9,]Z?ZdL-)XfNRQB5-K&)f<&.9?X#P?:BE09
1S@HUbQZVaD9ec^LCgF,X2F/+b+ZUK[>//<9a>LQbP#ATdVgPT4@/K6PDC7gB];N
)<8RN(Gf(EIH.NIK\&F=HFNG+Z<bG_(DZ)<WF4K5H-f_U]Sb5)BAeC:T_GS5_-FW
0-CD\7_bOO@/:TVV_ZO\Xa82JVX+V/9XH]VFC;JI7T:\@:0GK<P>FCBV-C8e4/..
I&;,WP#K,]dc2\[S9-82OcWL3,U;9Gcd3LD9[/WA]FKgS^.AO&Y#_-L3G)J+eb<+
T>NVIB/T#)#4Cb?(-_:#/)4R=F1SR:)PLC2=QKNXK&GdG.DR^P,HHK[Q8e_&E^96
Fd60;RNS[HVd^7)<_He]?Jf-0IP=^]2LfV4C1KURK#^R/4@J9ZW/D>B>LITV9aG#
?-9aY@KgBI\cVEJafU9:8M465gB&eI&[dC1UWQd6+D6_1RQ?D49?&5#)IK=W^@93
&ROd;\;9VBJ>>7G:#Xec.b;\I/8e>\:^:TE@Z;.d,XT/,[PGHIUO],-N(HXb]8Od
3IPdCVY+.F8ZP?_eBH();[M#AO:<V19CB<6<U&GBAQg2KXd=M+U+&?:=DT89=Z<U
\-=\7#FZ+;CAgYf>1&@+877Y[GBYJ6f+6gMO6W,]F3^Lg[@3)Z/@0:V:W3D(+=<[
.La6eg]85BIV71SK>&[4RfA1+@Y&E5S/.>RE=9g;aLN5TK45Y+9;<V5@e,Jd?AL4
#,)9R_;H]+bJ\[VQUUF;LG46[EP8&V/_5;b#:_W5GU2L:6&0C.@#a&^_P?0Af<(M
#W)eaTUGd=U5[9Y&AX6@3;;&AJ]A-];;9[9&@POJX.Pf4:129C4RE7VEeG=]/3KK
LHNVN;e),bLX9#V1]2#5S]3-4<=55X>OA;[?YM#gQWE\5_BcTXJNBacLc3ZQ+8RR
;<9MF4C&0\@4bU9K5T/f[BR):QY31#gLXX&WXJ)>)^MGe-L,dE+b-CB&dge9)X2\
DdgXK@e:I+^&12Bf97Z[0aA,[_SOBP.#&>L+fXa_W(g.YD1\1bZ\b-J<e@T8\dF_
OfKH.WVDGMSIEg70X2\.:S^L#R[I-427?X6<9BTBZ)WPEP9O,KJBJ8JC)f:?S.S=
A)DV]Aec_:1,&Z?gS2TX==.Ve1)cT0=P2RZV>M7?-C[TE^=]KdH6NXO/-YDgEN1G
[D,<8eb2DEQSRF^:Y348fD:&PXb=2BW)f<UUK&_:A[79GF6@8&F=KV_N\Ydfd6]Y
JPOWX][0EgZBEJAd.&A)/>f4,,#Hf9SH.Q0/eP#=d/[c_#9]aa>UJg,:8H&AORT6
L#6<)6@EKdfX3#8/QJ-F=/0fD[SN3+AVEd?<7gVfBfLbc29YRVNceT<>P24:?KC9
\>7+<MM#ALNR??Keabe^^^I5#)HU?[PNN3KOM1L#BP5JJ8S[d9=?beC3CLO<)YMf
3(-g0(d-(deGedNbIW<#&VNY7/=QX\.+7L5O52T8VZfd&(M&/A0EIbLFQ4&&:1,V
Y<@#)3WBLfH76?&LKbbEEbQ=[K/D>cK:QMU/P&\)[#>H^-Mc#K?QBSM,1V14)b-E
NcK1fg:cH5g/B83JM,K3C?f#[LW_2;&>(e4KE0Mf.DZ/2C7e;WERbPeYGF;OGW#_
fNe0>/;N#]52=a-eI3Wg.c_[_Y[A&XHZR;@Lg6JP:b7Xa9B&:FTTW51OV\:QV)G]
+H9/S])(4K&4KfGIS]LPNb\M8QH5]@P<-fV[#f_YD?_;R-Y<=c]W\C[6f,BI0680
9+R(DA5)R4C:)+dDE6=^T7F3FLIgVRB\eMUON0]cd+?EgU#X/g@L](K/#;=+AFB-
#ZbJ3BZIF7b<#RQ62,<KQXZ1DGUZ:G+U/.#Bgg<V#IUHEg25MHY1DG08QW@],WKA
,YMQQWDaY/+QF<JeHcQ+?_CUd#MJ,/8a#J^:@7L3dK_Z&dgd33e&&bG9<OYY<eZ#
Y/+4C(b#@0:e+)JZ5JXQ;?29gM-IFgKQ?Q;59LV/c&?RCV?^3=]JMOad^+<O7O=Z
,F&M(Gb[0eT&2[\:FOHV_.SN2U(1HU@Jb;e8AGXE;,6GcFGf?GG2+Gg+U6Tf?RE;
#EH7D/LDT5FTScKJGJUB\9>UHYM]1T?[G^.+P=X06</Tf/G/DD+T[(<WO6]H97M1
bE5Q7<OMDdEI4WXTCT?]f[]^:,GaA;7gDQ90-E4JC=7C6OSV5HP)OUW59=YB#^8A
,/:OcX(Y,:+e\YRDCUZ6NfSJc7BZf#eM>dH(\eG-2W#_NN\U7UgC?b+\8W1dbcW>
fA_@Vg)V>S<#C8PQKJ>U+TF^[:WeE0=WAPD,LaV:&4(W/PTNNeWS#Q8)X-CKR]F(
/O,2Z=aE<XPRJXLe-0aUJ@]>Ldd.A.aX0R3>#G&:fXIRff>?9G9YR-WAV/g,>R_E
M#BdB5MEX#21BS(+6dN3VGT(,PgR#U8,P;6GT,VTII?,3W_,e318YF]E8I++N+YO
#:G&/#TZV<#aGRAb8G&?-5H?g95A3eF:+)C>=e]]9X0<>B^T?/,g,DDcHGe0:/E8
\+b=dTNafVRJ0/d>J)NQ/]7A4FY1.GaCWV/Z1O=?+1C?[FM)M[MQ?,X.aMgC<XKU
G(eZI,CVf<2K&4.XK<bT9Q5[D:EDc>VZ\c5PR6<(6V/<DN[0G_CT?[_#8AAXc4af
L9dBT^H8=@Se^2gGF=Je2XZRK>2bG,H7@cM)GG@aLJ]>ef8:bTXVK.V[MfKL99_E
A:A5^B@e+\@gN_,2Q8/:ILD9IV3EL0HZBWTg/.2H0;Q?\VdX^G:HbY&LU[A0KG9&
FE<d1/L,4H0,10^Q-U::@@90fG4CU-CRgT/.HY<d2^T3VW[S<\6)VbL?J>gf=bAV
Ed0[UXB=G;/>\G@6X\?P@#588:L:IE4WY#O/Xb2bKA\/47a1CMM5&8TW](0IY2PL
(7f6=0aY.,f:11\GeIHDc7CK:0F21F(L_GbeRYOMDVEaZXTfW&Y80(DDF2gdfM>U
,>aIR.;?JY;:4+V9EW,KcD\5XI]+a0fgfAJ-\KRO7/3aDccSc;e)7ZW:JNaOYc-#
97Va6fKd#9,QeMBT:cN6<2UA?:D9Ja/;&fdC(J72;1>E&.?UM-=Q73/WU[TB(3JE
c7H2+4Y,,b(f#J;_L7#c-,52T7<,B?aJ#8YTO/]I6H]P:eN2K/[,:<a)KLM?R9#^
A3.ZCf:W5&>+&(7PX[\W646O8K\FT@<Q4HE]58-R=GBV?>[bU7.2P+JY[<?&_GP,
U&De7X)SAC\F<_CT>aX<BGJX5XP98:V6+^8>-VG<I(]#2ac1>DQe[9U8KdP+]C?<
SdGZ_\aJ])C_ECZ&L^)If7@^f3cb6&8XMX(aDFHGF:1&Ne6RT9HT++/[PROaV5a:
@4a.<^T2.;C>6?3V+@5EP-gRXCd((]?P3K;\&R/aM>J[aD1WS)X_&5eM_=DYgV<O
VVHa1-\NbEAK@FIaI)Q@54)7SY\MZ7_.R3ZE3;d@_W#[BE0NDT8B1Td[/fJY^X&4
RUV/3-(O;-Wa1(3Mb#Td&MP:ZI>VPFa+;444JS)SKOU-B4Q[\]_93gc+BSG\0,c\
fE/(]>EEY#E-)VaNGd7P#S;Sb@CM;H).&D^V)_g;ZJR<@aQe.Q0V^f)O66_.AINW
8ZXLZWN[D75;TgAW562&/CM;dJMGKE988TggOV&F9JC>g[EAeE9Y=+H<E,5L5X@8
bK#I-_/]A=Ab=0<P-ME.<W@320aC)ZUF@FeTY2\TdDUTVO^_bD7[b1AY18W8F50a
5>:BZACaN)cVfe2&)\ad:R9R96AHN?S])KF/6[-<ZM5We:Z13OK9K7<4M][XL/Mf
Xc0BCOQDb8.^?,g1D)GSN,fI<LDHPR^PR#B/O1_-KAH=,/W=fe:/,)5dCO>9^1-Y
A&b6,)@VG5b4/6RQKM>1Y-7:0W.GVVG3L<9b=MMEB,@3QAVLA[3:?LZaIM]IR@J[
\E5):2?DE6=P;\;6+/Cg]?f_-W</EP,JZS\L?gNTP#C8ECLJ2Q^^b^P:1E70,Dca
;4^^VdM.HDQ6GPAMR5)+ED/N,X>AG/HW_EMXAcgZc#CKUa/b0LNW(\0,0YFP(,6F
>Qa0(KP_Je2T\PW_fTY<7ELL<T8U^@02;+bB5>[M24KFEBcbGKS-F)O9&,ea_dBc
3H&L73QGT98&V(]]@;AT^X\EDN4V-&.B&-FC+2HX?c?ZJ2/Ge2.[Q);CPNe^fVQX
<>G4Y-af>2R#D>QA;.?)g\>D7V],)c6ab1C9?5V=>Q-]XZEF>dH4R#&<X_:Zfe[K
gbS(8VTPKXF3:eaA-+M0>JU6MV9M7MQf9cU=,)MgU0X0/Z4@)3;?9]E-V5^HGVag
d<?_a5FU5ZMHTNL@C>T69#/U+gg4#23&YYL-:GN6:&c=GeP=7MSg)bF=:c#^]#P[
58gVZ?N<U+&K[J3R#/.2(PYaP5b]-7WEIE./USSH1F=.W<,S3&W,G^:f]bY?;Cca
0&X#g0f831?PSPS7YX5aNFd3X8N<K:bC;N81B53Te8A).=9HIE\7L_A\A3fA;0eg
6_JI1^<]K2aO_T?ZR&)UC)FD(>aBN/LS4SE>fI+5SSSP<8g>M6&_@CR1HA;3T@Z[
KQJG]AA[+[bSY.K,\dGL\FGEN4&BFX?0\cO-M#COR5-NS:@@O/A1bZ64f3)e#3R.
.XeG4Q[G>4^d2W-#da?X?W.V8U81;+Zca8#2bX=:fLg)KP=VDNL,@QN=2)#HA(?8
Z>:4bW)+FgT]OUNH84L^15B_OSaPM<+4&3OBO-OF=6aK\?N_G5W2J6PIVX3)?Y5S
d8ZQ+Q1^_JDBF?RUENae@Z(fQ2PF.OG77A1E.Pg6KYe9C.\=;&0aIbM5_=.?;<X@
,&HH-X(eS7FCFU01a=PCf-CXC;@,=XE5X^W95F;a&934cdZ?Y[]T:D]^)a?/=[Ug
O#XYY=+UVfS.fc6V75E.f:f+B8T@f/89#J,@X8a8adU(WPMP?UE&?,^#eAH/58Rd
Y<?OQ+(:@OZ=PU+_fK0[6VHJPZ[(^f7_6&[^T\_@WD?M&[<6.BI[VYW?.6;T2RR;
3,cZ0QP2CN]H9O.(2B1\f9BJL7Q(BL7L;W3CC4AR@b>UcJdV+1A:H0[_R9fE295C
12?>5]/M+/=?c/1^)LG8:J.\;V]EaSXUGH[AQ>:&G.dTdQIJ-=,/LN:37,Rb<D>.
L]>SU,_f?8SR81-78<STSB+BY[EYdc)Q0B&-E<8YYZ\3c#+R]&&40];WO/b#2&<P
L)d&faZ640\f@_dJa5bB\=B8fe09,&dbS4G=-G>Yf7I?OIWfEKa=.DbYW3]1,<R-
GH)2#b2M5Q=7d?HT4P]Ug2Q56OGUN&]Pg?&VM(UI_7M9;d,;U+g?B9W-.-\gf/)&
?L?d75LD81=Q7ccX8[>(&/16#\@-H4CDXJ>JS)7T/ER6;2UG<<I2<3RN9:(#\[C9
)FTM5U4U5+LgRJ&Nc8>X1-3<1QW)YRFVT0>3]&dMC-A[+H??<7DFPESJXG[]BJe_
#HT\U+cLG325B2e_d5MAZZ87):ba>DV#2fX5B6XXfDT)aR_dLe+IePg#<feU8,D.
c(K3.@.)a,?2^7H,-BJbEMGf8[V?Y;WMHOBN.YUeD+Kg5cgf\b^(\<#KbL:Y>UJd
/R9CI0I+#QI=.\c82JCX4ad91dagL&U-]AGRHP1X[#FgHUMYaX@#]:U(R@Q@F5Mb
]F6e5LN2E6FaTR#,M@YF-T:)V\KKTAUKWSJ2HeK\@,]O]JLZa0:OM]bROYT#@M1c
GEQD:6YW?.E>RH:/IOKa19KWI^[C;+362A85:A1eZGFL0HRNgf-eTLfL1>)Y+GRT
.c<]ZCc,Y>a)+S4)Q/e[OA2C#^4DFQ)D782J#QJ9;dR^6U87(6EP1a;#B4E_0fZ>
2S<aSBg5D=31P?f>PN&7KUI;Lb>8MbS,DO1LHOfFR1PR(g=#]+3_7Cf7?2)d>(P/
_2d-;S.;/4_dEb7FO1_W4<9ITTS3-;=(82d<c(>I^Pc:Kf-.SKBcDP+SBVQ.f7V7
#TN/(_e]QU^QbO4e@f&M(::FP?#8<aPFXEV92Cb)Y46d#8MdI6e[J5]3[DB,O:NZ
8c0@_(ANFZ_O,5NC8gI(K_FCQVcJ2g5P7ZcQdOUY(X8U_>cFdYLCDTU]O(LEXe_#
O5:2@V#?-W_\2GA/X6X#+FT>;_J9&/[>71?2HZQ2L;1J+#-3?09&13_V[P(45IXe
.0G8e:FM0KLH>:8bNWFb2DNf\;_+3Ca0S@47VZB,HbW?XSA\.J-Pa65EB15C,eLY
5I<a^eKK_VdP&a3G>1DBO<,HSEH<^SSJb8GTF)OSS7VD+:6=GI);b9&?O0K,I9[#
;.SM<MX3T&O<eQK.FJ8bVd\F&6O^5O:(S#=Y,+A3()U#IMM>1+C^0U.H:2K1<NU@
d_>ABD:44Pf]->Y=bcCAMNS+(LHFFA;ULcMSIf5d6^KCePP/Z4b.<T^P+a@?]VHT
X8MB7G11.D^fdY/MfHUga7G?TfD>:^BS9[@.P<):=V>_(#DDSXJL[DA@IKeL8eFJ
/JCcWUc5\eS4[XcNOeS1Y(&2OUeHP#:P-Cd_0>&HDQEB3#&03NJH_1FG_?LSS&?G
+Y53K@]LV.)X[-0_HKD7:46bVeC3b@B##Ka,6PAJaQ=FA[U;&/?O7_+([JMF=[VJ
SW@aL.@NU1D<D\,4\#cH\[1HCT5YaKPL6HMWRO(JB_)1>V)/,1#Lf&^O@K?+f=SF
,R:b-97+JaMD8B<+F[7R^L[O<EXY(.c)0#eUT-6YbI-17P1U>Lb\GUHF)&JTCRLB
COY-STX2LKKdY,F+X,Z(e6Rd2T+3T@J[)e63EfN-G4gZ./C8YNG<2<M4LK>PN1+^
XZG#RC6bX=<0CDgQ[TYU6<VMAg]_,][IE6g1&7D[PLXaJ01?2=18^cZVTPga#H0G
S32C77DO/5&f?>?<HJG=1,aS69;1A<BNOaDJ#G8+K^&Kc7cKf?FI-^9aK<0.9_@9
CRAaZbTO0YV&BgUJLMO&,eF;@4f#\&&75LHa=1aBdf6D=M,6WT2GJ15J9<<0Q)/7
[)5OI_f]S-E;A,8,^G/=T^QZe0YL+7GA[Y5<5gXd<Q8JF_Y@3\Ta9g(&Hc=6\e?3
?>TNDO2B<D,)594^gY)Iea6bRY?L+ZLI43MdXO\?.Q#gG1W]U_LR#&C-X.F-S,HC
a(T^4CEcSG&Z\c_4IPYcS8R54C-#BSCFL:I=-=9,TJgKV\?/TZIaG6)[GXTN@^53
VIL5XRVcI[Zc5QYHHZ8Ge@03BcE+8O&b)^?MP4B4e];4EB7?/,7gb0]J4#<#XgCT
,VD#\[LME#+O=QQ+4I3^Lc_f;VNV9-070LR,]aMFbP\/a;Og=)\/F(cEOT^,.OWC
25Z7^A<bS:fMO6@3Y,8L#R@?Z:J5cF;:f;98XUVN5]<5d20#UAXY5a7.C5KQ5K-[
SR#?#4AQ(&8[eL.+SX<)&a[=>E=NZAVP_7[^=.LfS]331MB<9PH,YU.OP3AN0I\F
8EJ6O-^/#fYHE;dTQg3V-@+WEC@OcM5G;b9J2@-#2QZ\F\_O5/8=C0^M#QKZ14Of
@S<MfTFAH6K@R3#.,g]1UE4Ue>&5TZBEFD_.IT,^LSVSY,H-Y:]&f\cT;B<?0fQ+
U_Y1+?E>H.J(E-)[+>R<c0eZUQ+FW)cdS<dg1(>Zc4L\J#6W0F(-7LKL]=]ZUP2B
AIQ@a@>]L0b,.1QdFA^d-YaO6GG8O]LEBG_4gO16645ODSZ8/8]&ESQ=J]W_RBgR
g5MOF.CAVd;)2d727QX/Y1D/T\1?YA/4-Y?TC>CRDQ_?0:H;VZ/2e1KPL13c<:f]
\g5W9PK^,7I_X-?M<_7^gKYb-b\S<NPf\WUT(/44;]2GYIN><<^UI8OY6aNfG,S<
>04/G2bS1AffE(]H<,?Ne<MW[Z;(4eN]X5?EP7K:\@>Z5CZcYY:_]3MfCR\[fH=^
XT,dLTee?++-]W]&1[KbfQA@e/:_^/a.N?5NJ=A.6@)#0/d(#C;FJ+U<AH#HD+IN
;:&_eY;8&G328A8#+@UW,(JDKM\142J(,g.C5JaVV2&UI\:bJ0BH]4b]a8(+N(Zc
TH0,(--H_E[_TDNJWA;T8]0(<AQP[<7f7#+CD+I8NT/3)2F1I;U>5PdMC;N@(@GG
&IZ7d[03#19JM(:&\,</_HDO;>3d@5Ec//bgAd6+C6GG^dY3JZNbB#&XTC(gebR,
5H9Kc]=fWR.QX@I),3L]ER\RD<ADg80+(HQdKdIKcHRGZdS7P54R6J7Uc]F:ZSJR
B=/-SE2@eA;c-=JW0G/;),+O5VQ;4ATK:J&6KBX.RA/#cc\L+A8Z,DI/YW6,SW04
Y#UP=7RR=ANcU[cTaNdU5b],0=M.61USEc8-cdWBG.5,G+@ERL)E7OA,a;,#WJeH
WJE[9gcQXZ2(X]XP(/W:Kdc9d4)4^+HeQ3b1VV5Z1JREXGI_D]76+T.dIc,;Lgfb
Q7R/-I#-cCd^O;XT\Q,T@IN=eb;U8\g8eVBZZJ:D;)D(W&Oc7?=B36_#0MN+Q+FA
M)PVHbD+d,#c09&QC-F?DCE/]g^N6^0/U[)a+EcH)4@8CY=ZTM(Q/TGf(35H1f?G
UZ\>a;T#-?_;cd+V1A^F3.Ed=YT++O#Z[P>g[7dAB2?KTJ<Ff6gIBb9DNT5?M45D
X8Xd?DL2_gI]H_>><C-AcfNC]MBDKX_CCM0B6f;MI(d[?U\>,LJ@3LRb]NB_4A>e
IYPZBa0(#SbJ/d:+D[\--Z0_P4a<?@--J#Ig7Cf^@;NHJcD9O\?0)XB^J7,6<P]0
,9;^:CSMXc+Z>LIXfM7)YGX9PALC>GYEQ8(97H6<S57X&#+EH7D(\1@BbXH4]S;(
dP/bC)82a8AO3Y(Y?W.d7BcQ.00JO.SI/_eK#-EGgSNGDO\7#,XRTL(,3E5FM)DE
0[S]M4)FF07TD4[?5Dd:<B66UQWL[7?U;V?W9<Y)+;]WUO@ANcFF1Ra^eS)g;8<1
?^f6C/GXTRF)+R\Y1+a&_2?Hg96V8Z+HgGA:<XE.[A,[GXMDcfT)J][>^\_5>]QO
9]R=3WD4GD\Hd5E4^>+0._gB/];G<8C?IBYae=/^CKMPBAA(]I>>daT).]LM1gQ&
]_2[d29g[G909FZa3D\B:JZAUfdddY39#-Yb.R.D]bDK;;;LZG#d&X41)2#V,I=>
V;b&X(:F8^#UTFWdR,23W:[\aKa3U8dIOaB-YW];9;1c#Y/U7C=GgKZ;&a.;JW?b
_FK)2^6@@WYI3Q6c+W.YZHe(b&77,3-&8;ZLAOFZT@3D/bI1e-B<=Qe>+O]K:ZVV
eC5;a1+Q^1-LMH5-faWYS2IH1/O)ba6<b\Z)1/?e5VC4Zd@#PgJ&g&8S)5@]c=e_
N_bZ=5@:X\PWJE/Y[ff11R>V#V1A)D/cg62YXagOdT.NUa6]3D3TPR\UGI&]>I+M
SQZ.f+:,U)BZUHSZ2X25J##>>4H\^KJ@9c>Ge\9V1cTa7-XLD)VT2OV<;.U^N+gV
+bS44f]bM>c<Y5O&2GC<c#(>I;+@bK:-Sg8.(5=;7JW^=fK<9LW>>XUA\\b?LA&1
^UYgc3;EV<P6T18,Q0UO+SE.7L,=@TFaWND]&7YC[,^fY3__B)]NJY3Y0;c2A4W@
f.U-/f_2eU+DgLDg\N_9bNW^.]#)OJe\1\@.R#MV4DcVDOfUeX55,1=97&H-LF#?
4L3\g82+ZNBR\e:.2PNM(c4R^#/8,>g4<aa._-gZ68&9&?ES1(PGFN4;1T?Rd?OF
UbWVBg2VBD0GZ,S.2dcLcgY[cVfW+#F0Uc/H4L;N5Kd<^dSFZ:F1@aGccTZa+)4^
F,QF+e<HT0<<_45A4eOT7:F3b]:d4fG0b:&/9K1d0P7D<J1ec4)R-XF;LIMfG>aZ
40P02&4aY3RM>>VS?UcNcb@cLQ3\8XNH[9ZGMJPCP\#NcbU1bQ9c9;IGYM3]X6BE
O@)GCb697]=(:SG&=SQT:))::3GML]?H:<:_aUd9T@PZ^,.&Y3C\-U@:T\KaKQBK
,2g)@-43.1[>]=Y0@>5O9#M04H]GCR3NMaG]c/:=:Y8TK\KKS-N4UD#f7-dL[<Zf
-KFb5Z-D781>O^J4E4IddL-W[C(V/L0aZZ&aV0CL;X[+G3JZ8,U[M-:70_]ZeIAZ
88S5dX(T#/aVa9[K=2Dg6#fL8A.CX@ZK4IVS9.H[g^(=KDW;QW&-,g5]+LF(H;W.
cF4RSP@+=.D)>>fUI4H)ZdbIe0^V\UOYLQ.-;&Hc&MeL@GK+E[NAQggD71B@E_Jb
^)/IcJf+&,&@SK2#\BEYYCF8=f2UO]DbcVKYY?I,GZ#a?0VKV#9[Y(7[O<VKQG52
8^MUUSd.?S?1=X,S^ZX(NVSQJ-37OBI=X1QC2OIXKQ4M;.[C\ZB^:XE5QSQ]UFId
(0a/3Q^THcB=R0VB;K1@(AVO76B&GQ:6RFXVK8AYf<.^G2_EMM_8QD=]cP+@=TFU
&H6.)BT]U4KKF.eWQ;,S#Ae^>UV=)&MK>U0[=23bBG0[O]240(A\SN5_69)gTQ&X
_PO/Z:]?/+;g./MLcO>QGVH[5+O8PcJ^V>EMS;W7>aBaG/-K2fL/80^T.4\==Y6<
39]?cdCTC<58RZ8A27-S9<,6)aJ^O=2Ofb+/W&?H(T-A@N[6B,X61.c.W>7=]8D3
(gX:dHg=</+-A=,R2Q]FL420,Rb9W()>)U_.Q[+4Q,V6F\+F87^g18.Dc^0[EP.T
9/)+\MX0bP:>Q-S+fH>[NV?XF+&2#?WZDeXHV?Vbe+R-5W?[/413[,1f:-K\<7E=
,Ub,1c;gc#Zb:55:M(;8U(+Vd5T3G8C:208IUTF;d4E8S&V+^?#E=8575[N],ad)
NQX.c1A=L8Q2fWS_?6e5a<3eFeH)3\^fRa](Ce5>:,8d7SH>YNGbN0;33D1H_f/I
5gd+P<1F0fH-c+L&#3g8RM_H5QGd?4#<?<+U=VOT#H-YZYfW6SgAFNGfIP(U0<63
bB&L3Y91/1UP:&:eRN-#&)DES3f^(d6)SYRD1#\=dC95L/Y\CX6KE=:O&Qf_VCP9
M@H1)JZaf<B-]KYX+9G>D8ecYbKQ14YWXgUWCbTD8^WL^FSFNUI&FIWf?41H#aTf
RN_@25)JOB:Zg_J9W((@J\4K)3O5I[9E<cEJV6T66+bJT.,TY@)>F#-@&GHKGVX,
:1+SA;-4TS:][^X]gf5&QXXX2PSO>Q3a@L8,G@@ND.<>S3UgR9<7B07O.:I?Z9b@
OQg5S5eYKF/e]XH5B/U_c1cEWe7(\,=.[cK)=;VeRd3PQFE<-L\=IM8)VeCSJ4:C
,Ka76;H[(U(Z2(;9QV9RR_&dVd@bZ;S,Rf\b6083[B+@7]@Z#aBF(@T+M7OF8E@(
H_.CIGRUX&P?A&:[Odb57YOZ(_EOgb(>9>0:I?6(9\WO7?676(g_)Uc3CDW3O(;X
1Q=><#0^.XV03L?aPT]7T@0+IdR\XgZ:U,7Q0f]H]#Raa]EAM)UD]WP\NN2RC]aS
)cZ#&\VcIXO8g;EJT2g@+,KgZ>VbNe?MT1f6)=b4)/9K258R+L+edSUY1[Qf9]1C
=#H0D):Ma-R(eN4^>N<AZVGP/d5;9U?-I-.fA3EXM_<@T#YJ:)-aa>VVYKK6A+.]
N]bJg(:J9VX&HTgDYKZ<=5K6#-e@A9FV=g#//Kg3)3>765:S<6eSdB(EW(@Z9b(0
ZeMKV7)9PMR.AXaWPea-);Q<(c6-Q]aC1Ya5-L5:8#7-.P5J/&LP:JZ+f)3B(0/F
a^5X0Xe[M\:1FVEK=;\1BfUb3^A@5W@7J3O+D4Bd8+=QRVMQaI7U4ZM.e(N48>b^
;G(P=5TN)^J\HD]^=OKO[TJ),<E]./O:eO9/#1W?4VKO3>C]FFM.4,.1J20<8O_C
+<I9R5-6E0_[Z+3GGN+[\@Z7G/)HS7GMX1/1Y>cX\4\1fIA[>e[[:.ZC4T\[GA?R
>_Naa#\,5T/&dc-.4B[:BgU(=@;I1#YE@fL\UU,PA7@\D5+2e<0XAd.?U@;2M:7K
AY4DF,]=MSL;BP@PLb4A)&10BdE5AZ=[cf?RIL9f4E-A5&,b4WZTc]5_KgcTQ7V?
)D9&AaY/0:SF_A]R<E1YS6>[(aW_+NXRcO.F[MAK>0ZF=G:N<-/\:J?=4,TC\WaA
E[W-FGF88)CgS5X5MR>Y:QQQd8+,)->V/<Q4+A4H2IKHgYKe<=76GS[7\\+1<_TW
(=F8.5S695VNI8YM^G)G]_XAUB6=cJIM\KMV1,OH[:D)CX=/1Wd:)g@I0JKdXO@_
G9H3[.]Z5_4Y@L;,QW]bF4&5=b?/>+CVG5S5#BO]@SG_MeG8XU\E9(e]YQPSf+?2
I?Q&&_a.=2#Z\HK6a7@O&;>HF4>#XTXSQJXcVQc9^R1RIT=]?@c9-W-MaW?1C>b;
)^=GQ#D?SCU<-d;SbFRI:dG)--bYbg27@B][f:=aF=ge_+Hb]ZKAP8D5ET(I.PB0
837TOH)^F,(K<?+GfgD/2UYacYQ5>/MI-;.@@MM\4W?(f)c/eSf>0gZ-Vc#ee1RA
>a[g=-#R.R4RC2cZ?I-&b+F448=R,)ICL78f@L\g-f/HPagb[NE]J8]QEMbe):7;
[XeK5\)bJSWZaWP9857U/P81V^N+FO_#PT6?6C(W..V1:UcU8egIW;>NCQL:&/HN
F:e_3,JRCb/KcA@@TZ0Z##EH]]g2,=UfB2^Y\>5gI]HAA))K[,4E5b4@G.PGfPQL
/L\fA=EEA1E<361RQ7RKSc<4=N,]c4_Y;gE+-6X:V0FFP^XZG1\#@Id1PBcG<T1d
=L3O?SZY>ZgBU_F+ScM)[:==09#\COENFa6HH-CJF[^9gAdXI>H)AF=Vd6HWVGKY
D6,F-2#aKZ)9Y,(T3VB]fQ3-<EP2H)W]F?d</HR9JG@cWb;S:D72N@)>7YPA_NNf
+\VW(\>&Wd:AZ43(\Jbd3fA7aA4^SS_>[3QS/?-+9e_^:9]&;N^I5TBD1WEVW;#c
=G#VW]5]?SU&.=&P7#+_DJJCO)2DKSD&.J0W#7gWX622X[P.Q/=\g:;Ve7a4\0Af
Db0^VOf4WUc-6RG]Q?\BLaQN^L12>.USHDdRNc)-g5:(NR[H14G\I@3/M,:N:ReE
QQ0::[EA;AF0_R;=S>eHOMe^Z4_dYCFX[,SG3+aLPYFS@RKS/Gg,g&PP:aB_&K]>
E9D7IOCJOR0\5e^@1L1IY-La5L#aeP_;H#Y5)4OA,Z,_#5;c(OOe4Z-C6;S6ET_c
f3Y#g9(/+b0\#NER@f&[L9LL[ZJa14ee17fM+gY1BM/CFVY]0RAQD((20C3JAW0P
#GSFM@^L\MUK12KD^(Ee-VHT8)^7JH(UFa6ZNcSHN[DC:_9>aS]2<6\Ydb6+76=[
W90H^&M+S,7BBe,IC=VL&7c-PV@))b;2M:5Z?g8FAZGM0<=cN_(.O4.Tg-E97&C4
dRLNFY][d:J)Y0f,#)b1DTI3@Ob0^/dU9&DXM,&b2,O^PCRUgJ/aKGd.V-J=@H\I
e2CWgDE:M@A7AE6(f:bb1MYRFcET<dQ7#/ZJ,7Jc/(R>8_E:>NL8:M2P\68&J>ZS
?NB]H\]K4g=VEbbOT#9&YEHdg?^[Q350b7W?.0<IRZ2\SK-RK#7@D65dAR@N?_\1
_/2/72W3=CITT(QQ=34J?DAM9IU0XDY\#6_?90,b>>;72KBY0.;NB@B/LMN@EF6>
A6fBEEbM=#7dS.HAM,T@OUI/3^4Fe_Fb?)d]\]1[g/LXNKfUCDP7a[A6cAA;3[]I
aMHFR)7]D]0bJ^>gF>b,F(DgZ8&LKX^MYA=?e(=Y1PNA3K-U+]/HE9B[3.L]YU#@
ISbW32Q#Y8Z;bdV),>(O6L;NfT?P#85K>f0b?\J-?-<:2+P>@WX#[g(0AHHZZ.+#
HZV^NgAUgTA\WXA8\b6cO,=Re][ANd6[,H-MQ4MZdO?#OSeQ[-5^LJBK<=]WRgZf
P?[eKOKP[I&X<\ObMe1,-Y2CcVAQTe..<J=D(@=.7gC5;\1f#S_O[JcF7UU.b;E=
E<\(#WAcC<LST0S,G1YL_VWWAg76b#gdRKIM^\CDg_C4&:\EQ<O]VF^(58,ZE#+F
+0R2MgaI>cdPFH)3VOJP>&ZX&^1#RBE8[MWZFTD31-(3_e&dE=08+^TP]=9HX2QJ
cD?8F<C=<ZIFg1NPS-<NN^d^eE+^RCTf/(DTJKP;fVX(?E85.P-B-Z-#cX?M.9Q0
cHc&^RI,U0=^50(W2IaCWOD^L0MQM1+T?D^UG0S^1+f0TC)@:_4[CUJ-2&Cb.(d)
GDT-b9;;SK<_E.G)W3[1F5^_V3FZ#/QVcB14I6B]YbXDYYe;;5Oe[81>P[I.;[(6
@R,FV9^#1O?_]ST^7/0?5S[JOS/)8&73HW=8UM:].>aZ@B,FXW>f5@g7C,[HK,7.
CU@.XP#_f_Bf[72UZJ;33e8/3X,=D_,&Fe9LH<I<QQ\8b@a/A/RNATP#IM]_85Bg
g+S\X-308]C7Kg>^4/LYNOHEICI;P6NKX]\HG[V8<=TUV#]AERIg0:5cE7\XgWLa
cWLK9IO2D8<3^Q)?Y2\b\&7/+Oc;UU:bg[VEA.91V5F<?FE:@:Y?T1K]:_EH;e,;
a5E:=>51E#&:eB&.KZO5+\]JIZ4_^fRc69IH0O2^IO],R@G(:CEIJfVHR:2>MJ\N
F4-09e]&4KFBJ26O<T\N2J);6Mf\AAR4,+J_NR8T=IBdXI.Z?e7ZIN16-6S#I7RF
\S\-L7;KW\&&<I,CM[a].=IAA]#=Ta4U^fL(OH.Za1&Q>SU6(&)ONdbZ9)cDKA?Q
5N/;[4_F#XSMgZ5B/dB1#g8VI5/&;XF]Bc@OWJO(1QX>Q+-Y<(IG3E;ESE<)LE#Q
,JFHf,d6#:Uc/LY_)Z,4;53QV[]]#(LdKbT\(SJQG&D\.4:?,Y&LF[&FHVMKgAGT
0g7M+4G;)Gd7]:V0,89=<C+AKWNd[#1:/>U3S)b_+\T--2F<Z;G-.ICM64d?M?ee
;G?R,#@T58J=gJ#5,=1+27+GJF2=HF@>)\6F,JaUX502<.DJ[0NB?X1<+])4;,T^
9C8R:[(48e>9=1WM>N5d937dce^3HT.&#@<(TK:<YMIdB3E.I3=,NYZM^;e&JZ8)
Q5IW@6QYeKNgdK3;_+)T>1+Sae@Q=0A4f<d=c+OBJ=2;E5D>Bb9g^Ed]X5\Ef.Cb
M\Z[A9^.,WY3?a@65HWeH<V8,/QB.<QIKY1)2g<5P8;PKM5Db\CQ+d6Q?9<]TK\N
_M(<ULea.aP&Qg,1I,^OF1,]Q/D[Y&.YNeVMReb:9N1cVJAHX-^.6_?b]QSPE<_V
(S;71SG2:IXVRQ<3B4@_f?MdU4RR(Oa9=4O949-(;3KP+OV).ga^X18ZO,>M@6,F
US9,@V\P=E3TU,C&fS:Wc8J,0YT+]JP:-,;05VY9I[Q@A0,ecPfI0F2:0;ES\S[.
B7e;IeB(Rb/Ua[@6KT1cG/9[C0&GbYR#PB95O7_L_B\.c.FMHGL95K_aV9aAX33C
&STJbP)=ZY&XBPCNNI3cTMHe;0#6FM43K@afXgg<AU6a>510W^X7J&&)YGTIKL.#
ZVfWfJ?/AX9D=RA^>B;6[L03JH+VFU;TTZcB=0@ZF\896XCbB45A4N4Z<g6JP:S@
X1LZ47XVB;9[2W)&)CKFR4(JM]GMH(OBc7>DaYJ,L[FN?B^\7\ISQ4>-<>R]K9^;
6.Ia25>c1c1-QA0aT_QYf]P4]-YGT;_65UG\T8&P:#8L1H(3ReTb^>^[8]-48Rf+
F.Bc;7M,NFB3_^8XdN;F7Wa:T5_VI.__bC=Ye&H>#F(<d7>SZedVQV?fRacW8B6Q
(3fba[b=\\_Qf.?&:T.(=bc.?..U<XZ1[6H.4/.TI0#5:S9EX5Y?5\QA75YaQ]FH
D5ZN;2(Gd:+H-@IFVad3&2\Y-EW<EWf166QXP32N9)?S<c-G_G,VPL/#)D4WSRNY
gSI2124W92#]DXVU:ZA(01>0G]B7>cGG^E?M-A69Q)[LRR)Y1S)_K+>E=&7=@bdW
,D;[b2^LFeKaaK4=C6b)SXBRAbfdb]JD&(J@UF&2T>7?(#_)dbI\;=[6(bCH=dbf
PD)d_I0^8Z&g.X.M0XgR(HJT+98-)R6G)7dKBOFNARf@&)gP(.@ba3aM5O,aOgU^
XH5&V]P)HF5d.;6+>e,TVT[S@EYI;2gM&1bB>#/.-GbJ(@9aPc;2[7PKFJN--?V<
IN\G@X\<X_VTZ=11RDUFF>E6D#T9N(QP_^@Q-W4]94;1RdSbFP+5&T?.gg6;IH\-
1:O(FbUc<JMP;IRCKE6YUEfXN70+4_W,.JLd&,FL:<XbS.Ne#aD[_653HK:^I4-g
ZECIZS,KL<)+0ZK=(@D&OS6XC+>K_I\HIc=YLA3,=d,(O4)=]03](,Q+bO(1XbGc
IEa2NH7.g_ZZM?>@Ecb/P7&&8_H#:W>GJcP^+;.fZ0/SD?Ha>][AA\3)Fa.Vd#Y<
Z^YC]f]EGZZQ@S1LbO&dDA1:.#ZBFBY>XdR)/_d--d//8<I.YGL&5f+f3Yded]X6
)S\3ZI5aBWDS7N=1F.8;cB]SPBcRNOeZ:Q(JX[0PU25O[9cQb_6+-3W5Nd:(D<5-
?f^_?H^8#@W0BTe:/EI:14EbEebb7g6O14EOf.)39<=K2/YEgVS#,Z5RWB(^Xd<\
CfJ4WB:3d/TVVEWVJ-.<:Ge>c]-S^3&O)T6+FTF3d,UDg^T_+;fPL@JB-1/SA[V/
KH?X<>[8da+:d#Bb.HHfT_R-976/5-5@]0]4OK:O)7ER=RBZTM[X2N+]gg9bW;61
O7\DS,_)A;V[1-3d_fc#A3>07MG;+FC.[+c=CS6\<L<]/\=[>(X-ADX@R)NVAcO1
Z974?C.78BY+T9J94=(E/<O0PQLeZQVIc&8BWX_MB:2:RY4DeJ<@W0&?]5BXaC#X
LN^1Hd0FTLEaK6\5=3S&-.AW4FPDB)_/MF2SF6[L;QCSMH+3N-D?&bX-+&KPg9I7
?08:ff0?N@b,GR9^UZe?GWE3[H.5gNe+5/J18FFN_F5H]cB45M@/=F=+QbLXb4(G
MO)R#b(F=&-?642UGNRXeNQ2IKPUL4KJ9>d71+MIG:cfPL,Lc?P4(T<X+,.C(MM1
-g@HFF<?0@C@K5)fSBEHMMEXVHf;=S+D16L.g+ZKZa;AXD]L,S:#,=NODE^@;FFT
(3O<3BaOW/9Y_VH(bY[RGRcX_cMS+_(:-.1V)31[3FU>_/664b9FQ_](70@<)dM/
OE@GQ@6&G&T5U\\8U3aR4S;6:/FNMcd,0[W7NR6T?A-&:2MZQ4GLK0\7Q?3@fQZZ
5K[N;3;LIAC)a&Y>)Z<fZd4C#COGbF.2P<.4N2[^aEQ.>I;cK2&UL?OWf\dge..B
?+#eYI+;&H-L77>/OdL7TBW/WMXU&IY?NITJSe[Ub6,R8@^;0>H(_:_+DfSX7KB&
7Zd<C;3EXEHB)SM5<fT\_BCgQJHUC6.-)b1-H;9K?JBIb\L-0cP@IfLUM4_>978X
cd(]AI[B#3:?=)WD?dO\<SKPK)@/O=a_?g)G(D=J-^DBO6JdSCcfR?d]S?7-&1F9
cQ?UfbJY>I#RJBH_O?=>E\;B:J/)B(==[RV;c.SZ/#NE?JOR(U1Kf7eZ](1Y_&#_
7A1;)?EU(5dG]Ef7-:2)J2(6,eY-KWOT[dcYW#eM.5a;@#^PdW8-67Mb+V6?dg.:
D2J3YB4&RfdZN3([6E9f&5]F-P-(J,#J40V4,,J/FJ4_KAWYMX:>=Ce&a77,H9N/
K2G0WaW/;]3#9S1SK47>.Yd[E].A@d95JK#93Y>)_[b=X-cGMNLee?0IJe1;0VR]
_(affSL4L=TWB)SXG)ggA\Qf>3eeELR4,L0CH-<>,a4H,O.M1T78gADH3V#\+_9)
P:5=&-I;DQ\a]Sa?27AIId4??H+E4U9C7IA[O9O=G]LF86)C;?.U+7OBHNcYBT<6
J6Z0<9[W=N11:G3bIaM/;1cXA;DJ-3)[W@EVR(T8C56?AMDf;/1O4bG4Wcf=_L19
2H1gdC[Ed1F6D#N>Cd<Ia0BFO[Q?#TBV=gVRLKRf0^2M-7SLP69+=SO_+B9PfBTg
2f3_0SdO3?:b]>W)eU;&+20HKPGL]EGTKTWJX4:Gf4W#]_3</4C(2_G:Ob,2?KN@
1Y&IQCTT>g:\9OFgHL+237J?#3T#]DF#HAOYT;(Wf+NGQBL3S[K6>RD.7UbN/N\/
<-CQ9DN0>T,6F0?#-7R(#1;8&g279T)0=H4/XL>E;6fBL(D&,77c=EaWD_#?^e3=
0OMfeU_&Wf99E?B.7MM,^^3(==<C]QIXBXcG>;^H>?cM#dUd7+RDeP^O)cBBY;:)
Mf(,QME9&?/PW6;]I9bMHH]+,?J6g.-cGW5QYS3K3P8W5P0f/P6J>bF71];K4D\d
N[IQZ+2#+C>Qb<#E.C06]1O<e,>)eZ\<70^;g#M;JWHLQ.43\K-B71d=W7H(&M4O
6M^03S/,J?EU<,Df/E400](ETYXNCS,GD-GV?Z+-\R4feY_3,,BWH6:5D:c)B6OG
<UT5M,^P]BdO_9e5Je:H.VJFYf_-gSgL<5Wec>E+C-F<9Y<#AA;&@:eg8E^]&V2Y
2Z>(P,UG2?)CJf6@4JP8[Cb;D]f2,3dCA&_K0S#G5]O>XZ=OH3?JHU]JUc(JGM=3
8<V-.[38,bK74XF]bIY[d0=9#Ofe6YU/-W,aE:7)=F5QGD2=eD)#CV2UUE5-=I8S
DQ7XGcP3<?)Kf7\C-c7^L>7QP=TJA]+HV>B/dX+P)HM;TG;#_N=5ET<@,8A=+Jd0
bZC-+EYYUbOG9((L^Y0\>-QSL@=XKI8@f;QQ<OWG\DZ</7L\6?EICJ&?T+L553>F
Y]EZV_;AQ+S-,6BPSaL/ZbbgPKA9IPBC&eD#JJ6cT?]Ye[@AXP/+EeSY]AL)QGSS
FC@MV<\F,)#=HY;J5dOWT;FN/L:FR1g^&b6gY/&/I1,+2&\YB/JW5#\U.9N7^.8d
WMLe(IL7Ad2(ZW(8(Ug)1DeA0P,-QIJVMg6(#(/e&\6QL5Xc^OC7K6_/WEXQ1F),
.(aYA8.MKAG7BE/O.^5<5eT01V.+bG(B(CDZQ(+.^@PF)Q@(FXH4EO.1J\@]KSS4
S+^7PSeFPJL#ZfGC\:6;)JDC0EA^\GJTb@05AR1WKFR4Ib<FW3CD3.;fOR6D&4\;
7>PPI0YgKLJ[_7,##R2_Q&)&.9L(H16CS4#Kf^VNH<+3U9Q[#DTQ=F13G.XFL:;E
G,&\XB3eAZ+,PY0KL1RE)_EGd./,EZ(Q6RF,B)/_OK^((^R9UQ(X?@QgWMV^[FB5
a^Ld.)[WRPc1;6VS/TOJ+aI5]fV(06Z_QE:U4:UP=MHQ-X.f\0H.[Z^C:NL/M.dE
@b8ANeJ=WZ:1.4.Zf[+OR2NMa-_[_RMH,S^S5&7_W#Q(MGeX>d\1Ie;7_U\,YHB.
(#5U#RH_7BNQ&=cKYI>e7+a=4F9=E\#4,gb\G8WFVKM2KfF&\/3;f-Za2M1G?#CK
X1gfV:11/4FZ][If^L.MBF7-J2S&-3W0?+6?.?1>fAA4D_c.FcKWA?&^NY/-I+6_
341AXOf@H,@<2Z72IE\dH6<?(E]C\9D#\J+13)(Y9G8V[2V4U0[>?<NgD;R@33QJ
eUGL_WASS28CS_W;Y&R-11Nd[\1^03&XME01+X(CbRFDMO/T)AY\0T>0#B^,I+Ua
gO;9/5)WPd?Y>I)]-95TK2O7W7dDL21RgYOX(5VaD-b6Ae)e)X^?7-35e<&:\RIL
8g86_I=1\BI\:COVdMV\RR[R>\g;8-;&9D21AQfT^@W0]A/KJEb44HISbG--G0?A
8#6E;dW=<61daL<5R9U5&f)f&VBZ(TO2Z>#+6fGRJ#^J^)a\3AHd3CbN(_1R@<.9
OU)@.;3g<@\>0R+a#9[DCL-W8Gd6)N.PbH3RbgJPE3DZC2(80#]#e:X4LJ<7T.[[
)X,8cSXG8.UZAHL.1:>;aHBaa,(0G0/e8Y.EATEF]JU4f<:VIM0XXa^/ZPGX+L38
HP(7<V/JKb+aF2_:;K,WN)[FZ8-d&<b4@#3=UK5<1X>E88QH-Tb]+5e-]]R<d3H_
S@GAD>5AXQDW[\6XGb3<]U1aD/:.DPT+D-6KfL/aa5I/F.YXE#AOR28;7#7,0d/Q
H#N<,X(V<63IV8/S34)8?T\YN6dDJ)6-JJ6f7Q#F2b,?4b\B/ec5<Kc/)E6)T66U
0W2c7G+G[,=>_7G3ZJeQ+KgEcZ2V<YJT<W]S]1/D)DUU8fHEZ49&^6[(aB;M@KGc
:If:.QOMdA?J0-[H;[Y74[1Q/O5W>)0H2P3^FB=2gFM99Z1<XaL2<)b+2N>>PW.@
f3,]fB--A[/TZcB\bbIcU5)J/\AfYIPIXQ:4f(QZ8GX<b/_8\7fU[TGedc@f-L<g
fW?J<&I(SDObR>-e,(YUS#639,g08H^Q6+2.e[&6Ud3&^D@>\8gc);Tcd])TFG+=
3OK@Ed)7+1S.4T[afLV[[7=9]1/K&]S,8JaTOgI^#;e4[5QL8^AU+2?WYP7?:K<d
8R3CQYe#RSY6:G??WWe/Q:RID-LCaDcXK+1(-UM;1OQ\7/S1&8eg1P;9a3PH;IYZ
)OL78gR]Q3^E-#MUeT2g0R^Ce@Y;3S4P(40G[\b\3#F\YH7G+#F7,FRM.[R(.5/.
G.b(b^VHX-CX],7RAgPddd7ZWe+H7+3^HUIaEdS4dA\/W6MM1J-Ob254SL=Xa,bF
&^_dQ5S[+=6L<bg8GW=).]2JE:BfHb8V\2XMC>V5S-7N^Y8)VSXF-DP@KH#I(0dJ
-,d\,;YIJb::<G7:7(#Z;U@[L;^3c[EU\8Ag65Rg<YP++J@8@Q,^@Ka_A3AZ9=6S
dTc6.CN\IP;a[(.V><N[;f_JRGfWWX;9,Q(/EXcB@1.2R/IM.RS((e95&8RV?I7,
<f2P;Ag^,XT<;MFf.2D<OJb.4_^AeIHa&ISS17-:]GCKS)OVM3@2LZ?958<B1egC
IYDRNX^TOaG-<=8(e-:c<D)WV]<<X;9#YH-#ZLPN1YN#aU2XbH0fVK2>,Lbd7Y4_
>MK<OF_[R,BG2]O\Id@ccXB86CSWB805P.F.&GZe,X=dSf-D-DQ.b@C<FCR;8)g:
NKHc\WX1f;\H51LDT8aNf)70H^?54,+cbQcAU^Gd:ZZ(<N/4&ATEe0f&>/UF5K/P
XK;1+Gc&7;<@]A?ZG^1F@E[&+f(D5)Q](JK737:#AYMM8d,K;M4fB@NLC]>5+)TT
cDO:=QAf>6V70WO>8NN1M?I6)<d2O;SQ]c<H4-,;ZSX[e4f(ga&U;]CcNJKdO<-X
ECG+;7KNU#.3/dK>@B8LU7\[)CcP(N=30fXW)H.ZDB/#PL0IQBCJQ+XP2;-M0_?8
PIPDc4D;P=caV3c3B3&U[Pdgf:2[_AV0U0^\O/ag:-\7LCIcCR7g41]WXG8;,+_?
e&F>L^R^\K5LgOCIVO/:BDgD+K@KF?D^X<EaQ+ICTb12KA4?[#+U^6d\\(GT#Jgf
P8a_)1>M]aE03Y&6\)T#eK=O0@MF7M?d8TH/(_,V&)KbH#?.PQX#U2JYY<]b56HF
K;C/2QQ<af/LX:C=gMXDV[44>ASc4/I.UfU]a^aKf\F/^/dVQQU7.@a=CE^&Ue:9
.g6&Tb@W#1UUFD\,W=^8cE@H=CF,&_G\1Z_AC,2.96<UM8#B,c&C5eRb7-TQKdLI
6IKKRNZ&c]>]]FHd\()/,E3CKXFQ516b34XO=V)e;T.B:?FSQGJY,87M(V1+3Q77
2R#Pf^I/C3NL:ARK/3fC]I?M+QO<EFcW7&XfVR-X:I[+]egegK4O?].gY3+Df7U-
J^bfOR[cg?+Y)\a4)PRZ3L+0X@(N(f-_LSII4,S_^B@?(/g#H<QQ@>#VI+>\A:V4
]W,+e/1b^7K7C[:^B[M#CRZ[2Taf5X,;IL:)YV9ZOEUZJUee@?0Cc(H^S;PJ7H_&
2cBV_>b-gB&6cLd2/-VV0.BGTY\S@22FZAVfgCgAb\94X@),.,E<ZBJN^a>)FIeE
6Nd.L+0DUH<T)gK?^d?,)A4SHT+=/-94O?U-<DaEK+#1G/NJA?7F+2>/B.X[LM&#
T<:_4^VS5e5\<7cXdY)Pd9V1<S=]Z5Y3=d\3SINbb#)f+JQK[3613MHbXVdcS1I;
VXM)YR;0)FBbIT7>P,@0cI@;6U0#@TZD#EKacH76,LM[4^H2+2:3\<3UDbeG(I-J
0\Y/WRg(>f>Y^X@MA^LX\#5)O>#AK6gM6FAI=[95K3C-,@(_ZUa<&S2BQ]3be88W
&RK5JM3(M.3879Lf1--CeYC]FTRe(MT7H9fO=g(;&,+DN&Lb0IC/Fd:,JM:W^0b1
^fM1[FE#UL:@S1(?P[)I5HB5=+V=WKGf4X4fWO?V(cC]FZHW1^?C]0#:/.5gdTER
,X^D?b^SLIc<G0#M\TZSP^A?Z5SX;Q8S)3FHJLB&#UWRK.,0)I@YLLV\MU.LFMQ,
FIe/_@Ec)TbE:HM(g:DTD/cNA+P4H]=3HcPC</<=7;Y6Jd?W(0S@7aU&eUg7_03I
B2EV8UO30?TB+4eWPHLT[[V61]R.=0\NedH-]a^K&SM5+fb@-_1W3B&DCM7_]>)@
bR^fWZ;[Q=,P,f,^SA57Q09U>&(;#KX9,PFK,#bgO/WPd>+6Q-/E<V(,7-&e>U:E
JV716;E^G-Ld#SZ>P&.f6aLCO,Z@GJK9LKV5]OC>)=-Y6c4(@=&7CA7L>MWSZX:6
=U;J-:M4D25V8:fHES-;(9\7Zb=NUaC.@]\=+^>4,&NFVW@24/A+G@^NZ0<(TE#c
EDZ)UTV[W7?M/QEZ,];Ga:1VZ<XO<CE2NPgfAU9S.RHT&M9@L0HXfEW9EcK:[Qa>
)#>._\U<L]F/Mg7T.3^Z&f\F6^#395T:,0&[[<.1M81^cWLJV<U8-S00[\5]:.D2
1_#HT//^Z#D0(5R,XK[^Z_\-&D6&VM-58E&MAYG3P-B>M/T0bM@E:Y/W^<3L>4#^
=UWM;U(P9O<^/)_e[gfDNI?.Q]b\8Y[f<c?K8YROe8MZ7a6,a<;<,A.Y-/WUV&fK
aGCd^?7:PQMOL9,:2WG8PZ:2<]OQbD,Q)VfUKU\5&F37QQ/FM1[VCK9^F#efL-U=
fF>X1V3FbN(g2cC1H/UBM#0I>&NBGe7]f\/L@Icf6MPY60(F5ZW@16LS,0]@0fae
5:?\^60.3D.b<e))OaG#Q^/L.-HEV-DCW>L]Ia69XNP3S.EOGc8eP491W6-]Qc:5
NZ+1FWaGVH=7\E56#BZ4>VFJTMX>01_N7X6])VTTRPcEGGaE6S1-1XM;)X@S,IZ4
>-e,PL=gL[cYg[D7?^LM7Z5V^LNKJ,fcUM,Be]aF3C_54F[CL5_C20]EfNKH_NNL
8OA#K)/Q^.CRRe[-Z.[XF]4Sd_VJES]Z0IP.fb,>[UX\KgY:+@3GdXDM<=7\4bLb
1KO]X&JQZ7?M26_TcRMG1Y>e<T=;6@CV)(NVM]X@XEL(<:/ORA-c[=[([D@F9D+N
0]2]0Z.VB/K?LP.EI;^Y3]2M3ffDfA+2D_=E&W][A)dCKN]Sb(_#GX2gW\DgCGKB
cFOQ9(;_d4ZN,6bOe=FV^d;2#dfF..U0/#W#XcM?Q/fbJFD\TIZA4?=()(+=M/7;
0;f8(7[JY,8(F&.0H1\FYK_Ne3MRAaSB9HgL2ED?J^=a>-][>>B\DN46.N6:[T2>
(HWR2F7BT^M((8f\d6Vf\ICG1.4.5S;N/PZc-c?))6J[.5J_16QMG_0Fe]5,gTR9
60G:cTJa)Z\CNX1-PIc_Z;5Z1,G7K.._U[K,G:J(b#9OAKc#74FN=H^X)>2[XTDT
)&-&_KOZeVL7bOWUg9V/-CZb(K>8#PUF^X)?Z(8,DC,+O6DOSDeBKQQf>-#88a4J
)>59-QEYc&bOH7\8RG]>ZF(;fW2a<D>:g[UUQEERQ7V^MB^F1,LZ;-V(D4#RNcP_
FSc0c.ScENLY/B=;\GW)B+K@YVGYO.-HQ[:A8Q8^^&,-O0aKUF5EVLO^E2YC6++^
D;;WH8,@,O7Y1R8C)YFFLC##TAbb][\U6IITP#EcSX[OGTD0c&FW/=WaF0VY@55]
X40HOaQ/O=0VPKF3A<>=QVbETY9f?PC8TQ,b12@aQSDKgAJR0CEG_fY,XUA>3^FY
E.\g>;JDQI-Ma0U#^+7;PV^:3Lf&GHYRXHAC?=7#WOA]6A7[=46L[\R(&QaRY[5R
U.YBdJ?)IQJcGFHQMG7/7Y:P,,Gc2c,B=7>K<RMA;ON81:WfaCOHe)eVFR#8HN&X
-/=6?+GO.?^Y>ed<aFZ5&954a)F/;4V-FF]4T\[4f8RW6U[AO8(?a:d@+4;[=-K-
gH\)]&g_)[)C8;W#B>Q+9Ng/F+\U>K0;RP8GD5bM)XB>C4=Me=R&WEOGLY?=3>,:
d#&U(&bDU+0E[M^cM=IHV#SB<&6e,)g6R]EE9BM@7-M0&\M?8:.@X?5FNSO2b.TO
XCX8d5KOBC9^C6bSQd<5LB?3Hg1-N#(L[1#K=KU4<)4H5F3_-eW>/F.:KT,LEW[F
cE5,MIML-1VcUb(d8P7FT=+W#&AgG,23f#T&=OJ2JNb_F)Hg/T@1L[3#S(QJ2Kc@
4;_PNFR;W@GHbFCJ5#4?6V1S7>AC6EZN_F>SIF.:@KV06g>FLX6VSe:MccY+2_&g
MUcJ]H&V^Be;^=EFZT03H7]_d>\-JFV^V>6J5TNE>#d,@3A1Z:HH7A@fD&U.WXZW
<ZLP^[^c._7?d>N?H4WO]L=]1VMR35NQ@6\;f@^3>-55F\5GMU/Q/fMZ4U0\-QCQ
815Uf5.&&G??dXR7aVASFJSA+gf[KK4/QaLL+7HG+:EaQV,R716ac6-_S^>?VMdR
LTH->VEZPZ3d7J.BL<<05.6W]&/@SVTGX@ZDV5B)37)=5;8>B:/g4Z1GKJZHggXP
LU@@)6L?63_9=I-TTUVR3L=E&9HEC;W4Z0DVAHFY4J/UG8CRdBU/+4H5)JTESE#1
=3d>O_[+I]ab/?^;@]V@U-:OeR<f+6g)IG0>5RM2/DOJ;IVCH/T;+e[gLPe;O]aY
V5>-]M7fIUW<:MB;)S81/<>O\-,NV>7B4K5Tb=_76U^b6BYH]Ld_6?2O\-.);-,7
MM_D7)a_Tb72bRB8g9##UAE&f?NW8a<cQPR@+P:fT:@G#SLVeb;KDK)dgbJ(J=X=
O_[_;9?D1Ub@WHL8fSg+5M#OTSbO8AfZE#S-)>;UTU8I2YX(=fBT+:1#XM,=1&>S
KCNe/fC&:NYC0EN\/Y6D4gQ686A+>_Pb&O6(W9;(X[P1U0[S9&?ZFNUKcL]@953f
.J7ST)M1FN/:=0c#>[M<=U0P#ACKKPe=J7&@ae)[/NEF)\:d^)LJY=N>G>+fI&M[
M)b[B0Me^>/,/_;;EcUEKLTFPA_ND3O#K.5QgRS36cEMf0@^:A#a;F/bCY2&RX^9
bLEb&a/)6,b.-UO-[/QI?+A_c(G,S7)SXW(?.^E,DO7@ZcfYNNSX5+(OGFG<-/Ja
8Z[V/VHKSLJ-OZ?[@6:MgV6;G=.H+,_<9CHAZ1X^Q&e<AdHRS.X\V0A6[[@?Q2R[
2g-.eU/Q9:c/-7V,WRSP+G\15K=\bCLXXV7K)5DBK5Me1cD3d1A<OH2S=/S3<(cf
3Q0a[H-@ZYPPa&Q[AG:g#^(N4G;9E5fc8\[19,.>.Q;/Q4RVL2GTW&E;QJ)^L#(+
(?d4E41NS61@RW9Z,GF?CL8TU-Ve-+F]].f:O2Kd<<HDe7aP2N_J<#]XZF-G#T=<
K:b@\\INLIfAE4GW=].82#YS0ZS(Bf0<0O[?PVGZE@]H-]KQ<gEOWaR<\]+=&FEG
fbf?ZdfIZ-UJ+(SB=)B9e]G][==;Y/eL>2Y:d&UE_1\N?M0g6>58,FCVH+=&OYW#
RDSA@WY<#T^W8=N/Q9R81E<4O5aP28=\NJY6=fP;N\9LSN10a7-8Q)A)XYJ_/X\N
g4X,LG3]Xd1Z,92.+[E^Qb\R=dc2&+.G8UU<=H6Af\R=L,_<cg4IQNQ=\C>Vd6F[
7EN;d<g4-O4@BRDE#4PX171H]NC\_U_P+d&<0X@aeXQ@XRN>(=\]T<?3BR#1Ab8)
#BZCUC/#aeF2T73QQ2[a_\^(+)edY5=EK[HcbPCfZ+>b\e<=0K2VX1cVSgE]TLX^
]3)1LYU]]aP7S4I98B&fFDG[Gf_J,X\XN.=:c1e@_05[M[BI3S+^bfEB.9KZcE.9
J0^2SLBUP7ZTWUb_=T>d@T7T9<[C+J;JYgL_V377R8DVD8)3;GMZ=N(W_+Q^/UG2
@WfMB6SEZ5@U#STZRV0[=;f;E@D7P_FRdFB-@3/R_/]c,?f&XQ5Gd/?P>J5R)C)g
MHd;2d4e)Nd>X@e/XLHJEg-;dFP9cY1D7D[M5Q,)O(NA>fZ&Wg.G3c1[6>(8425/
T;R5a)?9VMWGS)2NMT[.>SG?)F\+UP.1V4)..HR_AY;9V]=KD#H8BQHcWa9>818N
DOgU2,50MJ#B)(D-BD/\S4]bFGa9cR&KHC2627dE#01B&14N2OM]HX2@d1a-->]Q
V(g1QVTN=da&P:RB.F1;;?&QNR3&PF@Z^OLO?S?SQH98S2ZSYF#4N.1a2f2d;)>g
N0g1@aP3[5S1CEQVO-@9&BWR,SWXALRN2?-QN)dKGVQIK:b6;+P0-f7;16XTd(]_
PIb/IaQJ[S25?GRfBPK<))4ZBG9eF67TV?<ZF:W#,;S-0Y4;Le+U9c45.VTLSU/8
TYF>Z\E+U1+XU=6]..\RWa9YC#7gdQIfL-3,a>3D6R?:^<8U^Y2Qe;&BQEDB>UfT
2SA9K4@I)fG7Z@KdE_P(,\aPD5ONJFG+.VNg+F/Me-W<[^)-^YCA9H\7d;7E9[@c
ST1VZIU6R\ZKI4EQMIc_<VXLgGP>5@M^>^U\,70A9T)g<R,Z.]C>(X__QP\U[\=;
5?GO<DF.J5Mc,(CUP.XRf]fN]<QOU&0\MRT0Z_D3IS<73OYTQaDH#dNVeMVQ,T?g
#0a6RdeW-QMNY+E1Z2/=6FBaDI1(>32MFN\Xb3JA6#7HPJ6O4E=QQ<RbTDRaEU[Y
L-Ubbb+5MbGY;FgV:<T_@L@I5CB9?e]708SV\A0/]K6FF\Mbb37AMHO>YLWR^8>W
=c-E5/;c1GEYB\a7U&V(Z+HRKJM[5.M>Q+7&4;:N\ZT4PJdH3Ya5g;W[#^^O&H/a
bP628]60;]S:QURWM0Z3Q]]A5Nf&S)A?IV95=^M1]+5BREGVX8KSO<Q2Y630U4_?
O3X:CL;@F;B;@E8D0GBWHL1N3[SRNG6(cAGHQUG(BHg[8O]W.U=,cXR[[/HgJ0,f
L2E^#X]9DKYe\I,B8964Z^TLB]1-5WYP8=)JMGR04Na,]1gF\fPW>g\N3K\9PY7_
F1&P.\1VU-BR)9aaa]6F29^]>ZY2:@ZdOeda88/Y=/RHQ?Lf#^L2cV(G:(WQ82@E
LYA86OSVcHUNaAbUL=^d/dCEbPUcR<>@XP0YXCSJV\FSO@RD-1g=KS4JU3;Cc@Z_
CPF8G)TBB.:)80^:TI6&8@fZ,NYP^bN,)9-.G5U8.I>eW?RFXRaWS<,ZJUZ+6YZ9
>/3T5J?..a\.Z4a+,?,?3]X3A1<Hd14\>+D6,0g<KR?QfN/VM0f1)\25&57?d1:H
^D36N]/67.2P4(O2#R:g;=>ZSF-EAU(UN0>7]d6XE79.BXB>cbT7T;&8_Y6D?MOB
[ScNaVOf,[bdBc8U0J0B0J4SD2#EUa)S.;8;@Y0f&K7c>(A5[_W]N6bg+,NLWb8E
T[b2)47&6R^@I?8XS57d3[1Q/34IP0O@cR(G(?bc>P87e-cWO0+20K][&,PaTP&7
_/+@bF:)(f_D?N,H0QC+R979)WWMMF99BGYGd-#?9456?b]W&d=C\SS-F9LC<V/G
2^581\#;>Rd_PZ>-=FM<BCZg8Z<_MP-aA+cceIf\eQPd9B/a3L(E;[OTcRN><=C4
e5/&/K]5X([+6bC]K6PDd/C67B?f[BWDMbf0=,_<IbLQ)X8Id:U3SP<_]T,:fYMJ
a,.15<f@/D5<J_(R&D8+7<8.:(:0g83G)VQ#J7#OAQ:WOKAUX--(:V1Kf(7F]>[U
K>a\+a4-Zg,(-XXa.LfY].5Q4IV^2Bg&&gXXEcJ<4:1UVC1.GFMME.<B4:[^-?NN
NegG:3@]WAF^[gPe.:b-Q9:@+]/AI+ISI-a;b]\7+PB4FJP=[T#A8PX8W]efGP:2
7aGB[UL5\fe&g5H[(Q5f9TA-7JGF3JH.Q7D=^X8UL]#\,SbV=DL,H2&0D_A]7>YO
.33U?J=6DRG/QNBDTf2?cB#)+/J8@)CI?M6.SX<Rg<]&R;Yf1A+,>UQ^9c/LB.G@
HWQ.eX)06]4E<)BCU0<^SUTAODANZKaV2\OL+Mg:)Ie,>FR4MR?NP;[2,..N(,L1
C2<Q=GDE(KcaF6b7QL\e3#F.)-/ZZe+.6^L&XY84RfgDV0C]ZXF[B=3d>DY2b=XY
E5JVQ(f/faNddPXGM@4a9Z^,]-L),1NC24HVfOI/>8J6K[bP9S<^I(TL@A=K=:UX
^M2;U(>L^(f1WPP7O\<?7E+_PB4\4Q:N/9?)UMGIAcB72bDV9\)JP6.d+8;LaG<L
<@TaQBP7=&P_RJ=WYRX\FMH7?9[5\6RTFBO/b?97\>eCgH,d:)1>DWaW<AJE3M5g
N0Q.ae:9Q07=PZD1F69=\e2d]<TV13H/_ZG_7L>bUa>b.G-;?DYO_H^)?>ZP+)1N
Sg5<01-cH7WFK4;(/TU,<T-b<)EBQagT;a_B8YbW&LKfV#X&/OHBU]1XZ8GgZ8OE
6(b,)3J+_#M]8B+Y3?Ha[WM#+Bf3D::3&<CGbaEQ#@.E6-;E3Y\+fQd,ed0QcQ^G
LfV]K2ZPd2RG@Zgd?7@:\9P>7NO=)f/Fd7Hf#]6\^DJ.46VL#D=G5=aS9@3G;6B-
XDJT#4N4e?\H<AIRO2F0,e<)V[7;<XBT;]NWTU;AEfA==4M-g+dZ:_+&5WFLV.S7
F5@_Y\ZNc3bZIFW,PRG9&dRXEaUJD9.#Te288(>W>40GEC3_faECM-dIfB?ELS[V
3V^8=;Y9Z82e:)(Q_1C67S+d:R9>RXaB3:W<O:EU^)?KF7IGKa18&M8O@4.W\7_P
+eYcf-Z4)cZ8c,UA48Ia)]YELb(Pb;_Z3LG6b5&Y1/Q;eJ=2XEZ/.b<U76BP]^35
=O\9_B^Z3[(-BP]M3^WLI94Z;UaePZ+c_T:LE#;<9,e(2YS:6XF_ZFSZ(WaVCZH(
+B#L;YL23QB]GS5\e7#QOW^a8e3[0#a8b;9TT9+&RU<Q/PX8e1>)Sd>fT44Qc6CE
F[3UOCW7bCT:X+4G]ceG3Q2?_C?##MSE^c&W>&7JeF-7]5]<[)SOB5R/,9Q2G8;3
G,g=H?)+cSPFT.T/(>ac^9.A2:[8LCJ<&T?O&\74@JK#3<Rf[5V_K,ZHc05O85.7
\FeO609=^5,^TL;XQEQL#3EW^80;QOG4CG]RWWN\\3TKC?N.R^-JeSa+Y[XG@=X3
Q<(#7(Ce]ebcd@<GCT#8DOT2;RC0V<JB1.)\,D2a[DJ5L(8HMXFG<T:.Z-aV>I1+
&E>g9]2JObHgF<(@V/R/.4FeMfGZ+ECT9>LKd7a]JH;#I8/^F5?:>GgAV96PO6E[
JPNR]BTfWQg)cVgdS9[Gd]b^B.(#S/1:6F:+65WC-5I.87HZPI;O-YMcCZ?F5<&)
a\58SEgb5.ASI_KKO30D6\Of7#65C&LSc9#Kb?8X7d3cH=SO5:6WJX9a=F3f\HVd
E\89fVK<c[@e+6R6EKOV(\XM?7eAeZ9?45[TGV29CWHGS1C8&>;?#g]W]Fd?LgMI
(aD^1ZAG.[?B4JQ=M)AP0:FY9)4V:LQH&O#EeE7-DfV6\@D(W>#D\M.50G/-g_e-
);[cR4Z5/J;Xd,b<g66F,GHX.0.5_SF:I=X7WKAb;=M2SV]gWT4=cPB7G8WKP\?c
47SJD^JaBDU7/2(_4:L4FDd2<;0WKbG?CZV7#)X@+O&6TJf8dY&S?LUZJ,OA&9PC
AgFd#:WT/]8.HSUQE7,ILG_I>#H3?Pe596Cb[gBVKaZe4UK)Y;M2cIA4AC##J0bJ
+CDLIMgb4\B.8&_U347_Qg7eDYDIZ\BW):W\Uce&X6A#TFAV)+]Q5M?TECRB[=_S
=1V6-P;<]fS.adWR@MaVPe9Z/>UZM5=-F_HI..E3TS[?T\0SdT=:/UDdV/NO2//M
3B>J/W_=..b824PLE)2FU=TfE4aUb&SgJ?_0RTPECM]P_^W2Y&dYZVXdKR+F3cST
D-KL<G(#K-EWY(_<I(g+dQ-W+^><=J41OOd0QIcUPG1VKd\@>+=7<gU1F#PEUb2@
5ED45T>-MN8c>Q0DIA#I.-T3,/4=bGM+\W0=R[MH4Xa#G(K+2/8[<BgNRW41Y\^#
#G4.>14V]U[@.cTV<>/e3O8aeO4R#ZK2X17&/WST&C,a-?Y\AH[SB>^A@3,>JdN8
ZNKB@:P#N\\OW+/6XD.)d5?W9PA+;?G?dB?(+W,E\6J6U<86@/UX7/B=<^F[GV-4
,=90Qa:edZf0C#+7&R0&e,2V:aUAWbNE@Cg7_=HXP^2,eGC)TbSaFTN@MdH^5:aG
I3+.VT1Q21-]2#F>2)(MMN96KQEXTc<IQDeGK6A:<S@gNZ+L+;&J6,gALaHR;4dX
eXgW/(5/D-;;+EH^eJ).9<7cd1-F=Af>,;9]/#b]Y(4CQGD3McIcJ=MA;a+HL)>3
NdO8EWM-aP(>_<X5e0P01\1)e]H1P44DG.UfFV2A4&9Bg81#9GcO:01^1O7;W^KJ
+/0bebV;E&IZS=V3QM=2H1#,>O=Y0RS0-2-/M##AfeAXgG0eS9RQX;LVPU?@G]9a
U]AY#QUDM@M&d9b()8QKg#N5f]X66@:@_#,,;b;Z@3^[V32\T/&Kb[[@dX.T?R8b
-c-c[-^W:9T+R_ENdcN<C38GbI;@8+8AWB#G66I=W#-#3,FeMd>T._Se?5C>dA.J
4I,>MMDA;)^OJVLV1b?8eB4M9>MVL#,5N&5LRLVg?D)?5=a5J8M\JZA<N6)4AVZ(
cM<O#_X?=F1D\NQ#a4^P?=983T,D]2KV2<T/_+9de8)<:P>7H\]\#E&,CIT])BI?
[_FV6FSB[+)#V\2Vb]-&&E=\ND>=T3deYX-a_L2)Q9KfbbWE]RL^KKB[NZ2<?_CC
30Q(1+5WSVW&T#T#,.WZeFR32K86d;:cLDA1ZPVP@>\L09:,e0UNB:Jd@.Y.+FHE
7C/]=72FB/4U^dF>9@NOH#^W3KN06ZD;eb1#<F^Rb>4FF#DV,(;;+Gg;)B2#YS/=
-62&c\_PR31#RBGAHQB7HLNBY<B[9JQKID4I[fZJWbb0b?A?Z0A.WKBYUN&[g9\/
9C6;\3WS.DAJRX(08O38E?Z\;+XTW3C)@e_F9eY.O4V5bG./YFg2@>2299;C5\>0
WgY:BE5\c,T=E(P]cZ(L(6cM2K:DH]JA5eIV]XOK&EQ/PR0)>3[W)IRJd\:U\9SR
ER#@S[Q2^.KfI=U0?K?ZK3V@KUcWC-&SQZH[[USbW[2e>R@=WS]WUX@+Q:HV<F2@
Z#e=-A69-bba2bDDK^eV)b4IWHcg6IH)Y2YQ5\]f[;a1>cMNa:.-RWH><d9&gaZ\
QIJRc6aK7f^S+gH1,O<HM\Y=A?_VN,[S2S0+4a)AdQEI?[:3JA;GYNXFKOM=5/MM
_\F<>P,F._<?=[c1Sbb81F.VGgE4e]HE8d_)OZ.(C-RI+eZ4VV<[[a&.T>JD@=81
/YY1\T.EZN_)1_?(S,JW^aPOe0(CX[^X>C_SDHFNH8[=D4<-_(dAbQW1JG:2XW)#
IV>F]F(6EN(9\(YMeP_ALW:V)D-D)Ng29BS>cJb7YMag+JI,,9.]0:&44fDV9C@:
M]AbIR05GY#L/_H_63Sd2c__#c&/>[<HB+52G;JQ9BD,:5^(gV[IZA7U0.RWRd/Z
B+BgF)H,JL:WP8LcZHRDS+XC+8/ZHV5UY5M@G?=bTb9[>f^5O_d[fHL8/4C<I(&7
.DQbcT-@HD+V=(:0\>6WaS;,H&C3+[7eQ7a#JE1].d5O#\U&PVcB1[:U?KL7)@3@
1.g#;3;CcJb>K=/e5KNCf>d94MILQL[_PFD-S&CIL6W8BB^&GS&^?:e?8E1F;2f(
5:=2_&5dMS@_1PC\Q(b&D><[O/-##]J35WOZWYE1LbUSbFVce;_BJ.X.95:Q;X_3
0V0dOOXZK(F>[=4bZbg+W81.((=R=40:8#9Df/L2<b)V<N7PI9\>U^=U^@7>1CLG
JE7T63-F?W1GLg6CW3b=bG0If83,2HXc.2O;GEK(cY<K98>_D\=S<IYFE[IGMCg#
GS0K+AH#,13HX)4?LE/5J5\P#(;WT8+D=5Y3HUdBDNcB[S5a0OX_KPVN3(,7AFgY
1a\;<dgE=Z>RaeGK83>;5P.e:bfYPgcQ>M607@@(0P1>D=U,U7K(-(68Ug\B1bQ=
7^7R5,)7[<#Jg;)32IIJU[ID70N759+<\HBVZP5K(a-L4.[fO@CQB0KOO,^c>a6P
+D0HQ;\fbd36gB.a=e\,[fDFZ\N[,P?U]I,>H^>=]N0-B<c#HJ]BS#\dW&L[<H,N
-R0gWXQDcNB&U#Wa#I4[]#7f,J((UF^[PM#f)dM8LTB;B?@<Y1)<O^6=EG.GSId?
;0S8d8L3e2-^g475Td\XO(?FeDLbEXL,AL1&&b2F5]?D?f\IV]X.V>[(dZ)]R_\J
HLF#T=7N[^E(1EF3Y@&Ma>#V\@,K41QYf:Y1X7:(&A8=R,ERWJ#@3@a1MY2;5eQO
AaL,cR=22:CZ]bZ##=Z@Pa_a:,6P3&TfNQ8(c^eCB957aJa[Db6773d[CN,RDZ0e
1SQ(=H#4Z20(eHHP-68NOdY.0C3_A&+9&.X+XC1,G6CL+:#9S:OSMecZ<2A06GaN
]cB09N:e^.]caANdb?E<_;L_27)59A9a14ET)&ODc5A725AVc3ON4]Lga^.d,]8V
Mb-dR=U2[T6)O(_d@1]M0GUgP1b1d:YgTSY#A>1Q[9M+)BGLC@FeU1Y&1LF^CWc[
/>7O&V&(^WG[[WHG8gCR1PHXM?K+M//1OW>T;4M_GA5VJ_2DPTL<U-d1BdMT[-F:
\:DI[G[AG3,9]L@(,g4UAS<W,TM@f#aC\-W,U&,]7b)fbCcBEc.J1Jcg.4#)+JeJ
<H=]C(L7eT^MTRb?YgP7/?\TaJ)&(N0Z.dMG:_8K=;fd@EYB)W(T04ZN=00\E?8U
6UWe\#YJ;6YZ^YN0&X_R^BIK+bHD==9GRc\51AQM+J@<#a4/Yb-#&+69T)07U+&&
8S3I^9>,SXXN9<A=QbdY8B/@(MF[DII-b)GaUF3>OU&HIL;6fg?0B/]P/SfY[838
5M[-bR#Tc;f=WU8OU[9e=539Bf2__fS0DRTBcX^X3T170BVdWE[H,cHZ==LWASP+
P7;V_M;7Na^4A+8J@KIccfU/NH-1RCLL]O#MYfV]7d,?9AJ<?&eb>\6TE0327eFF
I#f_QK^UK&5:5Y,R:IAQ/fA;#(#X2DVbR.//YBZTCBJ2[Yfda6SCVQ<NU1E4bF9Y
GYG5AJUbE,cO4(@C<\C4M/5e<5ITQA7EF?&0g?K_+SZ<<SA@/)K<+1Z]B5/(T400
]f2FJ)5F>IWd3N9,OBVB=#TV-D^<&bEPXdPe9bD95&NRdPEJ6cY?cJ\0ZW73#c>)
R<0=XHf[#^Jf2P6gdF4U<33I_]D<?>=HF<=PS&+ZOH=?MV/_##IPV-EG8O6:3]2/
KYKaJK4>aacXH7NN0GP+/MM=B[cdOTbZ&eM+bP72#EY.FVad-ZHbQ5;5D85WO@LG
BWdWH[,J9Z:-JQPA7AL34T?&.Ya;EF_,>Zc9=GXD4[LOL:PPN-D30([KQfGHM0:?
9QA:)[I)9D?WcXTb8-d/YY;+\)>=2BSgY8I2SaP8A9<OQG\KTLN>:&:D,;8XA0U(
>bFVP\?gMYK-;Md#1(-=#;Q0/5SAMGIX&1>Z<R@NP0c]X6dW;NSYMUVEfCL;JEW-
]F),D()1)#<]/C:UX49(?;O:GKYK+X]BQG\[SIN4/9[Q\T-YaD;0D0ZU+NNEDZ]U
M]D(PBN+)fW<PEPcQ5-2K@9])^[H)V/,)4V832Z)1GAV72^LGd:E]<=dfcVML#bc
/da-Qe,)]b)&(#)INWgR&?B>HK32PEdeRFXX.Qb,9OGfX1e4L0CN2-Ma)&fRKXJI
<HcHZGN:OZEBYT53@cN2I;Q0Dd&VcSf:OA:,ZM4?9AgYcRI>dFF5X+J+[?-M->SH
&85(LJ@T]]VgF^df;X<[PRD<X^25[fWLdE0<PQIBY?#[F2RU24@d??.XAR,e[Qc9
A\HA6:R)J[b]ZEYc&EEUQegS+g(E0#KdSGUW,0;F3VfTDRQB?ZD=@B(-4fA0.F,/
K[IKO]DZZHO1-@\M@U1G@:Z18a@bD]c/:10,#)QZVEFJ]927;38Z80O;RDHO_C;<
#0^DLPcY7Q,[/G\e,cf)\^5Ve&+(24,C3CF4AYb_U,d4eb):T.E>[<(a1IaeV>?B
_cQLT9#=ENVLP#+@)gMRT/fCIg#8E_&8^8ZMDLD4ff62WQF)G_MM]0c^V__7d<&A
57=V;Tc?ZN(dB3;ZBf<Y^OM?M=N3/T61>]\,1B.G<8(^XM13=e/FDCEDG^_IL,N+
K<KIX7980gUDP\NSa]Q.]EUL&YYZN<O83)V)e-fH>P,[KE__N9_AFOF5fT17g2\A
Y/G;-:V2?;c[eJdb?DQV+gcIW^)O-68bgE,>,9PVTL&FQgG>-9fb(B.4CNSGPB<_
(312YPIAFd&QFA>A<IKS4/:c9,XDSAZT5,_SgMX(19I?B-B?B^H.<MNA#K5=eRN+
L@<A;M_eJ]d36\:?X^=PAR5^FQ=;?<)Sga+3:M<,+V<Q.D\?F?cF8dS?;;5EEY(@
#9V-FfS>4(SObcV-,QYCD]>Q][?HP.8D5:FS;6G]g(D94GJ61PQPXL;K_;(gIE-U
W]BDH6ON&]J+1DC-BcKa,c17F2@W4GJMT]U\L?Hfb2a>/f=16(4T.gaGddR/8FLd
>-OgF-F>0M1D.XP<_fOZ[3UX?W[U&B+KMX)YP[NeCRQbUTH;T.T;)8G2HO)eHWG]
Kb-SG)FHFU)g\FUZ]QIQd^>gE>8,L&8XTE^JM>8CZT(JX)(8N-4@C/@P)P.?&<S\
(cDN#ccJU=;F3^:=E5:BJ&bX>^JP..-H09c@0YDOeA/S&8<#a2,&bHXX>Q;cBCd,
K0[P5-,Q_HKE^a>/daf;DK=YHF[R2+b6GgO;E?,RKHG7:0>MPB-7fK?:&W:E+FDV
T0_<W0C1HK:VA(C6I7M0U<5.HZf8\MZ.+M9-X5A&2,_O:/?1L#GZP\6-HY)DGKc^
7ME/g[/BB&5<fM\e?=BMY19Y[E(32TQSHIY1HV=G/59e6?a:=:G?.c<G2Z3Wd:=J
7R\A28bTT&dfL;[&P:6F\]>0Q1&<QR9(F0)AJ;&+P>Y2@5a;_1;1:H^-OR0.XgQ?
S4_2:_>&>JbgT&WReWP[.3g)S4c1YVOgVO/c/[:DgcE??[<8C_9F-D,U,IHYT/::
e=f\BM)Z&OX]=Q^?=^f@Mb.R+3(O/>&EAYBgI_F0MN5.BgS:8/6_..,C+642;b/5
fE+H4JG3>(3N\cQ_H/T3A/^C/4YF(]8#E92T_XQ=dB:\BD7BIEJ>=F3VeZYcMB8K
KKTBI_+ce+_&:/+^OROGJWT2W3EM9Bgb9ETGCBOUf?P?fD<F)7SLW4.Yd61[gVC?
IAc\(MD6FcM8Lc9V\I>3Y^TBTZ0C],JEKUHFaaK?]DA9cTY+Sa&]_DG8_L+GcR^_
cBeg5G0a-]S_+_HT.?L>?42ca<&JW:_.@2)PH-5BG;&18NTWT/LRG5--3@:L17VO
LWdBe+@#3Rb5/V@OPcbZ?P;aX[M(_;Pc^/:,=@EKe?-T#S?,0PgU7OG[?[fU/PDE
MgIW(HM+J@5T3:5f1&21.?A5]M?c@FX>cZ,(6fcPIE0e,:Q,TE[gW\0=W39J:R0]
T6d2\f>cPW:GDFYNg>66<><Q:5XBB:g=4\D\]QKV]#Y3F,De/QNIbG)@_@ZEWE,\
IJE@&O[6>9PZR-:dVZRXC-01d\7=FKT<g9fWW/]/eOG<?OPL_VODD#]XQ_b?7B&4
\e22HA-7GQfQ\QV&]Gf;UR6>>ZIHT:HFDe7P1(b&gT[_c(8E2Z[O[4P-0FfX-=1U
T,^[AM[LKYRc30,E5U;F6Ie0L)P?V7@6Jg5g:[bDUP?A#?5>aQM=U+_YEC3ROS2B
.EE6))d[,U^>AcE@JRF4gG7/P<Vc7LQA&5PB90>3a6[8\#R<^BF8PB9;:.2deZ8L
3Q1BNUOaGF\.63/Rd8[(<&=bHA_C;:&;B8/VV6b+Q[-,;f\+aBaOKJXBAW#SOI;N
\RY#ZPH^-9@<4>SO\1^O[<e>Bb1U\b;EJQQ>I(]:];RH<9_b[2(f#77D0Z<2cJ6J
H7+Q5H5>(19E?,X_Q0CKB@T3(G4029;KZQ.L/fWT\ag3:Fg.^cLAf@gK?>6[e=]J
AgOPAg[7:G<fGbW:_EXa7GE@KN(Q1?,0964ee=4d^&X,S?.cQBZ3V@]=67[<)B)L
4WJW>-Z&<I8C#WabU[bYSB8PPYg,CCU#Ld33W/]Ha-V^P-:;UeMN[T4FA=Y;1g4X
9A3JdTVLU2MRFAYgU]L,TbK&eS(/?14H[XA\]>CI>bI(]3W-8-XVC<_G#NF80YI.
VMaG[4\cWAbVDQZ+_97+P..20]W(BX<[4OCa#F.(HQ+-H0L#RE/]HO]X\&fRM@WT
1>P0O7]GS7JLbKF:U=-NgK<<1)UKV.;6(f)0]E-fbBXdg.QA\09T41-D<C5,^Q45
])6Cc0RD/=e2[dS>1XNgG8Y05?0I64]=((Aa4e/-:c[.SX0Y,eR7QRTLe&8U(>:[
#YO)2ZQ?ac,]0AIT9E:8[W4dQGc.(#:\aE:0F]H()L2I))0?fPOf-0aR:IIW.Z>?
1Tg3+UB9IZ_MS@^>efNFcBFc>@^X0;]P9OI<f)+95EfP_;@5(48/DU#G8Vbc(cZK
6UO<:?OCcbfcc)7AS]C+QX2[;N.[;?57O0(g9P>2e&P6SGALU9d>,CI(b(IAV-FI
TEVE,<+a1M,@Bd@MW/&&4H2^(dP9-FH>-5Tb>S/+NBN39^M5f5+M^_#[g5)Z6-QV
;E;(\HG-;7dQ(HQQ(H6cCXULH?BOb3BV6#JL_b,QM7U6R]P8#7O4.6)^QPIM2WdC
+J+)O1E\2/Dce4.,_1ZP5B@a?Vb>GLE5HTALfF8@WAa\Z].U\V4LV=Ae)MU?GJ;@
BMf_CQWJ@#XE+a6&Gg=a&&M:YOUec1CS0,CU&Vd/,=.M65cKH^ET=0/f>,KC4EI\
NOJGcL@QOWIf\)-^<B.g4OS,BX\OAN876N,QUYcZ3XJVRXWa09Fd_\CW8JI](R_?
7XVfL@OO&H&PfAY7J6DAW1W6O&CM5V+[[L8=88U[eeY4-ED0:1DMLeS0/J;R4f6Y
Q\GJ<34J8VPVF41BRW&O_NER1P9#8CHb4Ab_9Y+;N9R2b#3Z>Uce9/3\]fWT>2M^
;\A_]BB+GfAS#B41^C0edBF?/-d@TQ&3_#]/<.Q@R)>EM1Zd[X].M@D[X6;,Hc1[
X5>:Ta:+HSF?X^c4eDIZC>M:9M#UF&?Q9\?YK7?U2?ZEG$
`endprotected
