//ym
// // `include "../00_TESTBED/pseudo_DRAM.sv"
// `include "Usertype.sv"
// `define SEEDS 5487
// `define PAT_NUM_ 100000

// program automatic PATTERN(input clk, INF.PATTERN inf);
// import usertype::*;
// //================================================================
// // parameters & integer
// //================================================================
// parameter DRAM_p_r = "../00_TESTBED/DRAM/dram.dat";
// parameter MAX_CYCLE=1000;
// // parameter SEED = 7777;
// integer SEED = `SEEDS;
// // parameter PAT_NUM = 5400;
// integer PAT_NUM = `PAT_NUM_;
// integer pat = 0;
// integer index_check_num = 0;
// integer update_num = 0;
// integer check_valid_date_num = 0;
// integer latency = 0;
// integer total_latency = 0;
// reg[10*8:1] txt_green_prefix  = "\033[1;32m";
// reg[9*8:1]  reset_color       = "\033[1;0m";
// reg[10*8:1] txt_blue_prefix   = "\033[1;34m";
// //================================================================
// // wire & registers 
// //================================================================
// logic [7:0] golden_DRAM [((65536+8*256)-1):(65536+0)];  // 32 box
// Action act;
// Formula_Type formula;
// Mode mode;
// Month month;
// Day day;
// Data_No data_no;
// Warn_Msg warn_msg;

// Month dram_month;
// Day dram_day;


// logic [11:0] variations [0:3];
// logic [11:0] pattern_index [0:3];
// logic [11:0] dram_index [0:3];
// logic risk_warning_flag;
// logic date_warning_flag;
// logic data_warning_flag;
// //================================================================
// // class random
// //================================================================

// /**
//  * Class representing a random action.
//  */
// class random_act;
//     randc Action act_id;
//     constraint range{
//         act_id inside{Index_Check, Update, Check_Valid_Date};
//     }
// endclass



// class delay_random;
//     rand int delay;
//     function new (int seed);
//         this.srandom(seed);
//     endfunction
//     constraint limit{
//         delay inside{[0 : 3]};
//     }
// endclass

// delay_random delay_r = new(SEED);

// class random_date;
//     rand Month month;
//     rand Day day;
//     function new (seed);
//         this.srandom(seed);
//     endfunction

//     constraint limit{
//         month inside{[1 :12]};
//         if(month == 1 || month == 3 || month == 5 || month == 7 || month == 8 || month == 10 || month == 12)
//             day inside{[1 : 31]};
//         else if(month == 4 || month == 6 || month == 9 || month == 11)
//             day inside{[1 : 30]};
//         else
//             day inside{[1 : 28]};
//     }
// endclass

// random_date date_r = new(SEED);

// class random_data_no;
//     rand Data_No data_no;
//     function new (int seed);
//         this.srandom(seed);
//     endfunction
//     constraint limit{
//         data_no inside{[0 : 255]};
//     }
// endclass

// random_data_no data_no_r = new(SEED);

// class random_variations;
//     rand int variations;
//     function new (int seed);
//         this.srandom(seed);
//     endfunction
//     constraint limit{
//         variations inside{[0 : 4095]};
//     }
// endclass

// random_variations variations_r = new(SEED);






// initial begin
//     $readmemh(DRAM_p_r, golden_DRAM);
//     rst_task;
//     for(pat = 0; pat < PAT_NUM; pat++) begin
//         data_warning_flag = 0;
//         date_warning_flag = 0;
//         risk_warning_flag = 0;
//         Determine_Action;
//         case(act)
//             Index_Check:begin
//                 Input_Index_Check_task;
//             end
//             Update:begin
//                 Input_Update_task;
//             end
//             Check_Valid_Date:begin
//                 Input_Check_Valid_Date_task;
//             end
//         endcase
        
//         case(act)
//             Index_Check:begin
//                 Cal_Index_Check;
//             end
//             Update:begin
//                 Cal_Update_task;
//             end
//             Check_Valid_Date:begin
//                 Cal_Check_Valid_Date_task;
//             end
//         endcase
//         Wait_Output_Valid_task;
//         Check_Ans_task;
//         $display("%0sPASS PATTERN NO.%4d %0sCycles: %3d%0s",txt_blue_prefix, pat, txt_green_prefix, latency, reset_color);
//         @(negedge clk);
//     end
//     $display("============================================");
//     $display("              Congratulations               ");
//     $display("        You pass all the test cases!        ");
//     $display("        Total Latency: %d              ", total_latency);
//     $display("============================================");
//     // @(negedge clk);
//     $finish;
// end


// task Determine_Action;
//     if(pat >= 2700) begin
//         case(pat % 9)
//             // 0:act = Index_Check;
//             // 1:act = Index_Check;
//             // 2:act = Update;
//             // 3:act = Update;
//             // 4:act = Check_Valid_Date;
//             // 5:act = Check_Valid_Date;
//             // 6:act = Index_Check;
//             // 7:act = Check_Valid_Date;
//             // 8:act = Update;
//             8:act = Index_Check;
//             0:act = Index_Check;
//             1:act = Update;
//             2:act = Update;
//             3:act = Check_Valid_Date;
//             4:act = Check_Valid_Date;
//             5:act = Index_Check;
//             6:act = Check_Valid_Date;
//             7:act = Update;
//         endcase
//     end
//     else begin
//         act = Index_Check;
//     end
// endtask

// task Determine_Formula;
//     if(act == Index_Check) begin
//         case((index_check_num%24) / 3)
//             0:formula = Formula_A;
//             1:formula = Formula_B;
//             2:formula = Formula_C;
//             3:formula = Formula_D;
//             4:formula = Formula_E;
//             5:formula = Formula_F;
//             6:formula = Formula_G;
//             7:formula = Formula_H;
//         endcase
//     end
// endtask

// task Determine_Mode;
//     if(act == Index_Check) begin
//         case(index_check_num % 3)
//             0:mode = Insensitive;
//             1:mode = Normal;
//             2:mode = Sensitive;
//         endcase
//     end
// endtask

// task Wait_Output_Valid_task;
//     latency = 0;
//     while(inf.out_valid !== 1) begin
//         latency++;    
//         if(latency === MAX_CYCLE) begin
//             // $display("Wrong Answer");
//             $display("Latency >= 1000!!!!!!!!!!!");
//             // $finish;
//         end
//         @(negedge clk);
//     end
//     total_latency += latency;
// endtask

// task InValid_Delay;
//     delay_r.randomize();
//     repeat(0)@(negedge clk);
// endtask



// task Input_Index_Check_task;
//     Determine_Formula;
//     Determine_Mode;
//     inf.sel_action_valid = 1'b1;
//     inf.D.d_act[0] = act;
//     @(negedge clk);

//     inf.sel_action_valid = 1'b0;
//     inf.D.d_act[0] = 'dx;
//     InValid_Delay;
//     inf.formula_valid = 1'b1;
//     inf.D.d_formula[0] = formula;
//     @(negedge clk);

//     inf.formula_valid = 1'b0;
//     inf.D.d_formula[0] = 'dx;
//     InValid_Delay;
//     inf.mode_valid = 1'b1;
//     inf.D.d_mode[0] = mode;
//     @(negedge clk);

//     inf.mode_valid = 1'b0;
//     inf.D.d_mode[0] = 'dx;
//     InValid_Delay;
//     inf.date_valid = 1'b1;
//     date_r.randomize();
//     // if(pat<410) begin
//         inf.D.d_date[0] = {date_r.month, date_r.day};
//         {month, day} = {date_r.month, date_r.day};
//     // end
//     // else begin
//     //     inf.D.d_date[0] = {4'b0001, 5'b00001};
//     //     {month, day} = {4'b0001, 5'b00001};
//     // end
    
//     @(negedge clk);

//     inf.date_valid = 1'b0;
//     inf.D.d_date[0] = 'dx;
//     InValid_Delay;
//     inf.data_no_valid = 1'b1;
//     data_no_r.randomize();
//     inf.D.d_data_no[0] = data_no_r.data_no;
//     data_no = data_no_r.data_no;
//     @(negedge clk);

//     inf.data_no_valid = 1'b0;
//     inf.D.d_data_no[0] = 'dx;
//     InValid_Delay;
//     inf.index_valid = 1'b1;
//     variations_r.randomize();
//     inf.D.d_index[0] = variations_r.variations;
//     pattern_index[0] = variations_r.variations;
//     @(negedge clk);

//     inf.index_valid = 1'b0;
//     inf.D.d_data_no[0] = 'dx;
//     InValid_Delay;
//     inf.index_valid = 1'b1;
//     variations_r.randomize();
//     inf.D.d_index[0] = variations_r.variations;
//     pattern_index[1] = variations_r.variations;
//     @(negedge clk);

//     inf.index_valid = 1'b0;
//     inf.D.d_data_no[0] = 'dx;
//     InValid_Delay;
//     inf.index_valid = 1'b1;
//     variations_r.randomize();
//     inf.D.d_index[0] = variations_r.variations;
//     pattern_index[2] = variations_r.variations;
//     @(negedge clk);

//     inf.index_valid = 1'b0;
//     inf.D.d_data_no[0] = 'dx;
//     InValid_Delay;
//     inf.index_valid = 1'b1;
//     variations_r.randomize();
//     inf.D.d_index[0] = variations_r.variations;
//     pattern_index[3] = variations_r.variations;
//     @(negedge clk);

//     inf.index_valid = 1'b0;
//     index_check_num++;
// endtask

// task Input_Update_task;
//     inf.sel_action_valid = 1'b1;
//     inf.D.d_act[0] = act;
//     @(negedge clk);

//     inf.sel_action_valid = 1'b0;
//     inf.D.d_act[0] = 'dx;
//     InValid_Delay;
//     inf.date_valid = 1'b1;
//     date_r.randomize();
//     inf.D.d_date[0] = {date_r.month, date_r.day};
//     {month, day} = {date_r.month, date_r.day};
//     @(negedge clk);

//     inf.date_valid = 1'b0;
//     inf.D.d_date[0] = 'dx;
//     InValid_Delay;
//     inf.data_no_valid = 1'b1;
//     data_no_r.randomize();
//     inf.D.d_data_no[0] = data_no_r.data_no;
//     data_no = data_no_r.data_no;
//     @(negedge clk);

//     inf.data_no_valid = 1'b0;
//     inf.D.d_data_no[0] = 'dx;
//     InValid_Delay;
//     inf.index_valid = 1'b1;
//     variations_r.randomize();
//     inf.D.d_index[0] = variations_r.variations;
//     variations[0] = variations_r.variations;
//     @(negedge clk);

//     inf.index_valid = 1'b0;
//     InValid_Delay;
//     inf.D.d_index[0] = 'dx;
//     inf.index_valid = 1'b1;
//     variations_r.randomize();
//     inf.D.d_index[0] = variations_r.variations;
//     variations[1] = variations_r.variations;
//     @(negedge clk);

//     inf.index_valid = 1'b0;
//     inf.D.d_index[0] = 'dx;
//     InValid_Delay;
//     inf.index_valid = 1'b1;
//     variations_r.randomize();
//     inf.D.d_index[0] = variations_r.variations;
//     variations[2] = variations_r.variations;
//     @(negedge clk);

//     inf.index_valid = 1'b0;
//     inf.D.d_index[0] = 'dx;
//     InValid_Delay;
//     inf.index_valid = 1'b1;
//     variations_r.randomize();
//     inf.D.d_index[0] = variations_r.variations;
//     variations[3] = variations_r.variations;
//     @(negedge clk);

//     inf.index_valid = 1'b0;
//     inf.D.d_index[0] = 'dx;
//     update_num++;
// endtask

// task Input_Check_Valid_Date_task;
//     inf.sel_action_valid = 1'b1;
//     inf.D.d_act[0] = act;
//     @(negedge clk);

//     inf.sel_action_valid = 1'b0;
//     inf.D.d_act[0] = 'dx;
//     InValid_Delay;
//     inf.date_valid = 1'b1;
//     date_r.randomize();
//     inf.D.d_date[0] = {date_r.month, date_r.day};
//     {month, day} = {date_r.month, date_r.day};
//     @(negedge clk);

//     inf.date_valid = 1'b0;
//     inf.D.d_date[0] = 'dx;
//     InValid_Delay;
//     inf.data_no_valid = 1'b1;
//     data_no_r.randomize();
//     inf.D.d_data_no[0] = data_no_r.data_no;
//     data_no = data_no_r.data_no;
//     @(negedge clk);

//     inf.data_no_valid = 1'b0;
//     check_valid_date_num++;
// endtask

// // task Get_dram_data;
// assign dram_day = golden_DRAM[17'h10000 + (8*data_no)];
// assign dram_index[3] = {golden_DRAM[17'h10000 + (8*data_no) + 2][3:0], golden_DRAM[17'h10000 + (8*data_no) + 1]};
// assign dram_index[2] = {golden_DRAM[17'h10000 + (8*data_no) + 3], golden_DRAM[17'h10000 + (8*data_no) + 2][7:4]};
// assign dram_month    = golden_DRAM[17'h10000 + (8*data_no) + 4];
// assign dram_index[1] = {golden_DRAM[17'h10000 + (8*data_no) + 6][3:0], golden_DRAM[17'h10000 + (8*data_no) + 5]};
// assign dram_index[0] = {golden_DRAM[17'h10000 + (8*data_no) + 7], golden_DRAM[17'h10000 + (8*data_no) + 6][7:4]};
// // endtask

// logic [13:0] R;
// logic [11:0] dram_sort_result [0:3];
// logic [11:0] G [0:3];
// logic [11:0] G_sort_result [0:3];

// assign G[0] = (dram_index[0] >= pattern_index[0]) ? (dram_index[0] - pattern_index[0]) : (pattern_index[0] - dram_index[0]);
// assign G[1] = (dram_index[1] >= pattern_index[1]) ? (dram_index[1] - pattern_index[1]) : (pattern_index[1] - dram_index[1]);
// assign G[2] = (dram_index[2] >= pattern_index[2]) ? (dram_index[2] - pattern_index[2]) : (pattern_index[2] - dram_index[2]);
// assign G[3] = (dram_index[3] >= pattern_index[3]) ? (dram_index[3] - pattern_index[3]) : (pattern_index[3] - dram_index[3]);


// // SORT4_MAX_and_MIN I(.in0(dram_index[0]), .in1(dram_index[1]), .in2(dram_index[2]), .in3(dram_index[3]), .out0(dram_sort_result[0]), .out1(dram_sort_result[1]), .out2(dram_sort_result[2]), .out3(dram_sort_result[3]));
// // SORT4_MAX_and_MIN G(.in0(G[0]), .in1(G[1]), .in2(G[2]), .in3(G[3]), .out0(G_sort_result[0]), .out1(G_sort_result[1]), .out2(G_sort_result[2]), .out3(G_sort_result[3]));

// assign {dram_sort_result[0], dram_sort_result[1], dram_sort_result[2], dram_sort_result[3]} = sort_max_min(dram_index[0], dram_index[1], dram_index[2], dram_index[3]);
// assign {G_sort_result[0], G_sort_result[1], G_sort_result[2], G_sort_result[3]} = sort_max_min(G[0], G[1], G[2], G[3]);


// logic [11:0] threadhold;




// task Determine_Threadhold;
//     threadhold = 0;
//     case(formula)
//         Formula_A, Formula_C: begin
//             case(mode)
//                 Insensitive: threadhold = 2047;
//                 Normal: threadhold = 1023;
//                 Sensitive: threadhold = 511;
//             endcase
//         end
//         Formula_B: begin
//             case(mode)
//                 Insensitive: threadhold = 800;
//                 Normal: threadhold = 400;
//                 Sensitive: threadhold = 200;
//             endcase
//         end
//         Formula_D, Formula_E: begin
//             case(mode)
//                 Insensitive: threadhold = 3;
//                 Normal: threadhold = 2;
//                 Sensitive: threadhold = 1;
//             endcase
//         end
//         Formula_F, Formula_G, Formula_H: begin
//             case(mode)
//                 Insensitive: threadhold = 800;
//                 Normal: threadhold = 400;
//                 Sensitive: threadhold = 200;
//             endcase
//         end
//     endcase
// endtask

// task Cal_Index_Check;
    
//     case(formula)
//         Formula_A:begin
//             R = (dram_index[0] + dram_index[1] + dram_index[2] + dram_index[3]) / 4;
//         end
//         Formula_B:begin
//            R = dram_sort_result[0] - dram_sort_result[3];
//         end 
//         Formula_D:begin
//             R = (dram_index[0] >= 2047) + (dram_index[1] >= 2047) + (dram_index[2] >= 2047) + (dram_index[3] >= 2047);
//         end
//         Formula_C:begin
//             R = dram_sort_result[3];
//         end
//         Formula_E:begin
//             R = (dram_index[0] >= pattern_index[0]) + (dram_index[1] >= pattern_index[1]) + (dram_index[2] >= pattern_index[2]) + (dram_index[3] >= pattern_index[3]);
//         end
//         Formula_F:begin
//             R = (G_sort_result[1] + G_sort_result[2] + G_sort_result[3]) / 3;
//         end
//         Formula_G:begin
//             R = (G_sort_result[3] / 2) + (G_sort_result[2] / 4) + (G_sort_result[1] / 4);
//         end
//         Formula_H:begin
//             R = (G[0] + G[1] + G[2] + G[3]) / 4;
//         end
//     endcase

//     Determine_Threadhold;           

//     if(R >= threadhold) begin
//         risk_warning_flag = 1;
//     end
//     else begin
//         risk_warning_flag = 0;
//     end

//     if(month < dram_month || (month == dram_month && day < dram_day)) begin
//         date_warning_flag = 1;
//     end
//     else begin
//         date_warning_flag = 0;
//     end
// endtask

// task Cal_Check_Valid_Date_task;
//     if(month < dram_month || (month == dram_month && day < dram_day)) begin
//         date_warning_flag = 1;
//     end
//     else begin
//         date_warning_flag = 0;
//     end
// endtask

// logic [12:0] update_result [0:3];
// logic [11:0] write_back_index [0:3];
// task Cal_Update_task;


//     update_result[0] = {1'b0, dram_index[0]} + {variations[0][11], variations[0]};
//     update_result[1] = {1'b0, dram_index[1]} + {variations[1][11], variations[1]};
//     update_result[2] = {1'b0, dram_index[2]} + {variations[2][11], variations[2]};
//     update_result[3] = {1'b0, dram_index[3]} + {variations[3][11], variations[3]};

//     write_back_index[0] = (update_result[0][12]) ? (variations[0][11] ? 0 : 4095) : update_result[0][11:0];
//     write_back_index[1] = (update_result[1][12]) ? (variations[1][11] ? 0 : 4095) : update_result[1][11:0];
//     write_back_index[2] = (update_result[2][12]) ? (variations[2][11] ? 0 : 4095) : update_result[2][11:0];
//     write_back_index[3] = (update_result[3][12]) ? (variations[3][11] ? 0 : 4095) : update_result[3][11:0];

//     data_warning_flag = (update_result[0][12] | update_result[1][12] | update_result[2][12] | update_result[3][12]) ? 1 : 0;

//     //write back to dram
//     golden_DRAM[17'h10000 + (8*data_no)] = day;
//     {golden_DRAM[17'h10000 + (8*data_no) + 2][3:0], golden_DRAM[17'h10000 + (8*data_no) + 1]} = write_back_index[3];
//     {golden_DRAM[17'h10000 + (8*data_no) + 3], golden_DRAM[17'h10000 + (8*data_no) + 2][7:4]} = write_back_index[2];
//     golden_DRAM[17'h10000 + (8*data_no) + 4] = month;
//     {golden_DRAM[17'h10000 + (8*data_no) + 6][3:0], golden_DRAM[17'h10000 + (8*data_no) + 5]} = write_back_index[1];
//     {golden_DRAM[17'h10000 + (8*data_no) + 7], golden_DRAM[17'h10000 + (8*data_no) + 6][7:4]} = write_back_index[0];


// endtask







// task Check_Ans_task;
//     case(act)
//         Index_Check:begin
//             if(date_warning_flag === 1 && (inf.warn_msg !==Date_Warn || inf.complete !== 0)) begin
//                 $display("Wrong Answer");
//                 $display("Date_Warn_Index_Check");
//                 $finish;
//             end
//             else if((risk_warning_flag === 1 && date_warning_flag !== 1) && (inf.warn_msg !==Risk_Warn || inf.complete !== 0)) begin
//                 $display("Wrong Answer");
//                 $display("Risk_Warn_Index_Check");
//                 $finish;
//             end
//             else if((risk_warning_flag === 0 && date_warning_flag === 0) && (inf.warn_msg !== No_Warn || inf.complete !== 1)) begin
//                 $display("Wrong Answer");
//                 $display("No_Warn_Index_Check");
//                 $display("formula: %d", formula);
//                 $display("mode: %d", mode);
//                 $finish;
//             end
//         end
//         Update:begin
//             if((data_warning_flag === 1) && (inf.warn_msg !== Data_Warn || inf.complete !== 0)) begin
//                 $display("Wrong Answer");
//                 $display("Update_Data_Warn");
//                 $finish;
//             end
//             else if((data_warning_flag === 0 )&&(inf.warn_msg !== No_Warn || inf.complete !== 1)) begin
//                 $display("Wrong Answer");
//                 $display("Update_No_Warn");
//                 $finish;
//             end
//         end
//         Check_Valid_Date:begin
//             if(date_warning_flag === 1 && (inf.warn_msg !== Date_Warn || inf.complete !== 0)) begin
//                 $display("Wrong Answer");
//                 $display("Date_Warn_Check_Valid_Date");
//                 $finish;
//             end
//             else if((date_warning_flag === 0) &&(inf.warn_msg !== No_Warn || inf.complete !== 1)) begin
//                 $display("Wrong Answer");
//                 $display("No_Warn_Check_Valid_Date");
//                 $finish;
//             end
//         end
//     endcase


// endtask











// task rst_task;
//     inf.rst_n = 1'b1;
//     inf.sel_action_valid = 1'b0;
//     inf.formula_valid = 1'b0;
//     inf.mode_valid = 1'b0;
//     inf.date_valid = 1'b0;
//     inf.data_no_valid = 1'b0;
//     inf.index_valid = 1'b0;
//     inf.D = 'bx;
    
//     #1;
//     inf.rst_n = 1'b0;
//     #(15);
//     inf.rst_n = 1'b1;
//     #1;
//     if(inf.out_valid !== 0 || inf.warn_msg !== 0 || inf.complete !== 0) begin
//         $display("Wrong Answer");
//         $display("RST");
//         $finish;
//     end
//     repeat(1)@(negedge clk);
// endtask





// function [47:0] sort_max_min;
//     input [11:0] in0, in1, in2, in3;

//     logic [11:0] max,max00, max01,max02, max03, mid0,mid1, min, min00, min01, min02, min03;
//     begin
//         max00 = in0 >= in1 ? in0 : in1;
//         min00 = in0 >= in1 ? in1 : in0;
//         max01 = in2 >= in3 ? in2 : in3;
//         min01 = in2 >= in3 ? in3 : in2;

//         max = max00 >= max01 ? max00 : max01;
//         mid0 = max00 >= max01 ? max01 : max00;
//         min = min00 >= min01 ? min01 : min00;
//         mid1 = min00 >= min01 ? min00 : min01;

//         sort_max_min = {max, mid0, mid1, min};
//     end
    
// endfunction













// endprogram



//ph

// // `include "../00_TESTBED/pseudo_DRAM.sv"
// `include "Usertype.sv"

// `define TOTAL_PATNUM  50000
// `define SEEDS 9527
// `define cycle_time 3.4

// program automatic PATTERN(input clk, INF.PATTERN inf);

// `protected
// BG6QF\3O<H=I^8SJ_57UH<#-4&_ea9GeKWUc(@PM]b#B>X\19[ZM-)Q-(:^;=f22
// B&e_Q7Qc)FO=A3YU.Z]1XI5(OI>[eFDO=#b=O)YNOHFCRG@2PWRNJP0[TQ=/cZC]
// /9:AUA4>Db965E-cLE11\[)d_4#U5YQ&U&+],Q-;T+f&H?A3KTO[)X..S0ANBbWV
// fJN.]:Q4=I5,D7Gfd9QdCAG^?-FT3Jg_8\M=1/b9=KY?Ma0AO3BZ.3N&VK4#OcOb
// :6+Sf/OBA:6Bg_23O7VV0HTc5_-cSIC(]FLU[e8B/T0bgU(@XW3GeR/PfUaW)(IT
// (DWd\5V?/ZS\C(:TXH0<H=?.?+\O;QPB,Xf(T)OAd>W6Q7BJTFZO40FX26\M^&Gb
// (gM48D(W(cLUF<fT7(K,e3[+b)8OXVL(<33?CIfN3g5_KcP34;H?fGK4NG/DG0(J
// M)M6]dMa1(;bF0Ga3R][.R\K\=XG(W=Y3F=\Y:IQD3/Tg.DT3HLa]LMGIF@5G_5O
// )K;;;O^=:>]<]L=@A??7XM2:d1^\P?;0b&;bOV?&#N.gY#C.F9^b:#DV0EFSR766
// X=3&?>BH6\T,OBXF<KBGI9MH7(N=K<]&+NC.7M:+>df_O\[V4+]:TY0ERYF#1=3H
// 77[NaYT3MS^,KN2NA7ZBMaH<7(<UfTdT?Je]=LV](EF9NV>4(\@&LAQSc89FZ/R.
// GEd:-V2W)>ZT69\+=^-:N6_\Sf>6?,:-<<\U(ge5eRO^=::MF[ceL7_K2D0-)FB;
// >R(13=UOaG4L)GR0Fc53(]R#^I]F36d;RN]Ue&X53F=L+ff<7@f+UK-EO:2/Xb#^
// aIc;4C<AW0Gg4b<(=NL4M5-eZ)cFNaI9[=9g=>6>?BW@/&:=B9B\4.,LEB=eEDd^
// +/Db3-g5T1.HULRH4R<S/88=g#:)W4c[M\N\_FF8c9-Cda>Ka[8\Y1^1-,8ULdP=
// ;PR6-B\f6T/\M[0W?#NVUQ=??f1(GP<=@L-M^fX(BAa2V>VCKLGYM=Y++5L[SO&P
// J^GM2BNN0MH?3I\RV48&6@;@#,a5>da1=OFUT#ONW;UDdOL(6\e3->\Kf6S7T5&W
// :gPD?:D)2YN=egJ\]FAaGI88gY?K<Wc#]4@+C[5.QYHVRS@\LM.6P)A>IB[2KQ8Z
// [_0FMbdAWXAg=J8DX]a>ZRd:0J=1VBP-7:](]2V7FLG2gQe7)/:_6R9(@50<]5^2
// [@GJGZX7WE#[I3Y<aAc-IU4U1G/@.\THPeX:26If;=<78Q9YRFDG.Nfg5XQ;3B6E
// 3d:f7Y23#=g:RKZJDG;a_0-I3gIE?2[H2>#ePPZ+-YbX^;+/9O82EV/a\Y)3-ZL[
// c3&d,8X^\@^PMAEVF5^8Cb],3)Y8>Lb?HB(V62bU9CEIGYDQ1e[O(C#Dg-X+T)g.
// ML5AWK/<CFa,G_)JfTJM=AFA(P#+]Lc1Be6E1fWOWV9>B[+#5=I1g:Zg2W2D6<N1
// g<F2XdYN159dLNEGc:C9Qca9C;M^NMaT>6gYL4_TH+ZZ\_PeO3aWc]eKPA=1CO\1
// RBMI]>AQ)X491cC9,Ae)W8X?&f6W-?(U+[XX7AN81WUZ\Uf]&D7VG4Ag:+,PN[:S
// PLcU5#?CGYJU_;OJU^@507):<X:(JfL@[P5EWB(O&Y4)^b61^cU&eU@SOQ5>fS=X
// ^J-?Na,Z[I#;6JFIO3@g>#7ZQU:WE0BIZ=4e?JVTPG/<#(XO:&:cA/#[(3^UQ+,W
// ]LMD7T@cA-D@7Qc5\Hd?4cGY)B37gYa2Q4^TSU8SJcT#9Y]QA.d5fSOYaeNV;Ig8
// NU>CPIXW7\6@Hgc:+@I92-R2M+M_(9_<dW4CMDgESfO^.-Dg2]<BU72?A_)HV(OX
// 5cN+34Md(L:;HJP>)b#L0=/Uc&fYNRHUBT)=/UYWb/aB0X\?a^<>:?SZ?6RIeBVX
// 69\1WFA2QJ4E+cV[=S^QdQ_>\IID.c_+3,;+9dMSI\AK.[9d?FT_8X^2gg9MLZ&>
// VGgCN8_P^R^3M2?U[QY7(_TM0g@B\DW7b>fB8\#Yg.5=AD8(QMX]/Ha5CO(1./-V
// If@1Vf_<,NU^QOPLPb=7Q0?&6Uf?M\a9-0\JdeJA>XWUM[;2Lf49?HG8,]fWHUXL
// #>&T9a#S+32]8))J+5KBT/-Q>Jb+H^+O2M(]d,N\J1W^L^L&9::3>FEUATfGRI<X
// ]S-R,];_cA3=,@[5OXQ4d:I)M&4S<OVf8\#;S2S#dY.cE154EU^gFTd?<;0QDQa^
// 4]QOQFF+/23&fOI]34XN(VO>8SP0A#QB6(L:>Z,c1SX/23[fEQ(KSSL(fE.5;D&/
// We+FXCAI@-H&G8(5ET:23/M3ZW@I.?^U-USU3?#G=-TOQZ4Ya))NUQR?Yg2C=[UK
// JV98.:ITHg&H,:/#=3dPcRKP(K.N-/4L8Xe_;D3?@a(W30IZ>=cHEH0-TEI]WT4P
// RD,:[[-A>dd<5)FC6[F(BZ=6F:?O:216Dg+U6dA4d(3ET1,e&,?.Q3LH\RPZ9A#?
// Y]N_DZ-e].PIJ4QR?77-7-X[W6XY7g;f(Z-UAA,IJ9Q2V+BOf7K7bVb.f:L7^0g)
// ;3M\ATT#=6dZFK90bDOL]=DgJCI(L<SV<a+A>QbOL0U:HBE..+5M.B8AU\b2.gVX
// >INVO1YKEf[g34^KGUYcS;W++S96.2Ba1TETf6d,<HG+R2&e1J5WcKN#(YaL7_3]
// KQ;XDgO\dODX;+Gc3VReb,WY,FG,Y&d)9#WXWQ&&M4CJeYS+4eeEP=b?+#6bNSKc
// H>a)/]QXP03KU([HAf+^P0_89S)-Yg5RWOgQ)W3M.81F;;JV\=QD_@Z8ZB+9]ZS&
// EXWD\7f53]\8#[RE-M/25\RbVJ4\-dc:]@YPOS(>:TZ8L)=F-EP3QL2a(O#FDCF<
// =ET0W6]KfR#,@Vb2G<6&bK,/?@ddQ(XST8BD,b/1=CY6ee9bL^7,Ug1UcT?;JE[<
// ;P5]YES:<VD:a@_6U&).HS<&PHOQAbB)42M4>fC@5-fGbN?VNB((]WgDX_N1[KM1
// VGM9g-6?:gKI=]QOa)X]2Q9<]4&eb68>^&HLeWL?.KA4/5K?]6:H[5B7B@a^S9YB
// GY#/C8GODE>dX2].Y8K[eUSBNe5Z>M^e\XXXRUQ-INL9d6S#ACA.(K7H[;17F,QW
// 9Lg8I.X+b-R6#Qa1(S1aK]dP9e41d^/+I^I7FX0BEJa]-Q(;MCSPQb7<[B2eC8U-
// J\6>J<fHC=XD5R2)^_L/NL[c(DO4BC-9L-XReH4bYQ=9\P9/;B=eO/<f[bP<=MWL
// VgQY(]9^JL;J[NYZ#/.AS52Xe,0fbfJC,EGY^g&6bIAd#Pf-MfK^F>0e4S/.<I^G
// f18KR=:O.IARd;KXdJaOU)N&X<(MH.dDX#[XB\X#JLUL;)c08#a@HM^]^#U9,(+:
// Q>B)86^C\AUZHY,^e2>,(c-5635d<QKN8\8_N7_-VP8gKE[cN;f@]YL;bP+0_JMA
// @>dG(/V3FU)C3BJ_I-]R61>#F@>f1@P<@<PB+Pec2CO[O()b)SNcAfZ:7Sg:6SR1
// W9:<eNUdgA.b8YSEP6N<Z7?:3#eg&X(J7.S7-1gFU>I<P2C_2+_HEL\gXYR)bR-A
// _4VOQ-@T@cGK8LY)+Y2/7gO#2<7(GO83?&2=6fXdL4+SWAc)2^17<XTU[GT7N<O:
// +eBHfbE?L4=^Q^HT,Z->ccSR2LbZ@K4.&:4;QGc2/Q8<1R3Tf1[)0&C=O6SZ).bE
// L]Pa31EdOgK3gH)Q]RLYKS;A2PCMMCY7_-Tad(J[.g;cLVX1#U<UJ=Q-VDKUTf+f
// EX3N=ED]H)aJaPS4;-;gB(Y</W.Tc59IZC:;9?^CXc+9E7/+VVMg#.2.M85V2DR6
// F&7YJ6eF-c_Rg:cQ08E<S)OBI7,fM^ce.=DS_8Ce\WFMZ[2bR6VT9]\Gb#5JU4JK
// TO5MQAZOOU<3S^_108:c;2b7_AcWX\6/2C9GIF5>-W(,<6X26,(GbM5?aeQ.M_10
// dEB59>3fFB5c)TT)G=@S=]eC3#bU2C_RT1:P#7SCHL9@2HPQ2H&b7aE4<47CIaH-
// N:H(L/A07F@Kc7dIb##3Q6PVbPa3C#OY[G3A(<e8ceFZgUS::93ePS]I.R@IJV11
// )_./L-R?6CAV=OP+:TQZXe6G=;c(@9U+G(8=OR?_#P33]A.FgaYZ(F2B0>(LU8&J
// 4Q2GB.W&2_7RI\]Q>A0E\QXKUe44LH^&BaO8EKH.:8f/:FO=bWXXF=E+6YNJ@@DO
// C9H8LN_#/KWIV>IcaKX3gBc0&I#&DZ32#,)2V,J?LcacZU-KU:Y@cG-G=S(b0+XH
// NQFa7eQQ#EeJC98f>12aJT8)Jg1E&(eXE8VbBCPXfVd4\N]G0fc11dUd3H,GR3CQ
// c](Ff/dI0bJ82N;&6299QZENE)DEEE_+aP;+Re/c6M>H\PP//8N\7cWF3#L\0+-P
// Td;^FRH7GJT\W/I7?2@9L7.RR7Qd4\54@B;L7WL?34bHdGMcX1Oc+g)57QdW]gO1
// &b0&9aQ42:(IH9Id\XH@(]9FS/Ia7ULLCWZRNe9g]:6:aL=X/Rg(f71+:W.PD.34
// XWZ@=Pd@M:-[8&C,K^LBR_JRFf2SU^Sd/f.-P;H@N9e=BMg+7)4I<]ZEaUg7CeET
// f4;Z9g6\^E6#=F,VaScFJ0W3V;_3ZJ(F-RN>Xg7Y]\_)WLS:aHgdWDRfZaJf?/f9
// V:4M(SP50.@1M);g1#]c\EG.gF]U9=7ADG,UZ46R11f9E,7;5;UC]WE?MH=6R1GR
// JDc^&)W5RfB5=EW<WCJ43W<eTPa^E#B1RH4D^cP?21#7SA]]OB@5d2N:TGUJPZ_E
// @MB<\L7>]+Q&:<gJ6<>9bA+LaZJR+O4a24\8\OT<TY[)O[+<VT<)[M)L9JAUc;IA
// 5\[F(^LK_3DK7>=d_e256Z=U<1K3^0V+P@cDg+Z)#O_1-^G&?92)g2XSGc8=T0[3
// 4R#VAT)Bc01SZF.T3]/<XNA5S>,22U@f7U8AP>]2P+CD24EU;R^:F[#),dX-&<T2
// VD\ZCXcQ2_YJGO5Y)Z<B8IW9CL9>@1,&;)C1;L:>c=PFeTY]F9GU7Y/(0M:8E5==
// I7Da)VA)Z9e4.6\F(R51/Bf2M]/aQ47E7V3.VfSCFM3KU(/V+_>+AK)4&&JCQ4X;
// 647.B^LfX+beIP>ZgX/ZY#5EHI@G2_8L[VFSR>N]C57,-E^UL<@Q;TfJ^^3BLBGL
// <&\-/#YO^g;&U#<COYX>]H2^UQbV1ebOR[D[.#D]V&CeHD?b.].KH?e/<S\V-WKQ
// C2Ib;XLT?1D9OFE>N;W]PREQD142QSR[M0F_AG2DGH)I;QZXJ/_[D5OaRFRA1=]K
// ddaFaQL>,;C?TZ;6U@RLCe][aU&>>&A#9W2].,MD(JX(0&10<PL1/OJ_G=_Yb0Qa
// (D6[-+?RAE3effU02O<MP.+9H5G]6Og9Z^DNR9.@aHK0cKZbN&L-_[JD#-LD2GX_
// 9EAIO^R9&f[9>HdW1T)0@=@T.G_FeIbE)gQ\P@JMKSA:Y9&?890<,O6,0dJ0)QcO
// (SE7#c(>WXN]b?2^)43K\>M;@J3>ZRA9C0HTbgPHe56^d\<NN:HL6Fb<b93U+@YT
// bfSIa\[;YdW/K8E28X2Ic(.=c4WTN_@KVH/Q#O5#2K4e+@eOK);B4S=3#P30(<8)
// Wd?5+\JF&Ue\JW/N=3GZ3E=7>cb+ROM\FA#W4E>eAZUG^#=?8U)#bR>[R]CEU5B7
// 6Hd13Q3H3YOFO&463YKE101U_@5>X&&^f??&VV^^#Ue[a?R\[L[/7#ZCTEX#(I4T
// CHd?=W]J)->-Z.]F-@(N]/=Wa2V6M:&\.Z:;5AZRI>&OOO>>Y84D,M\_[Z/9eV4L
// )DX448S+H;_>Qfe6/f1(\);c<&T;4O+9Z64YeO,^-N>]#9.HfRgR>05=R]@@.-JG
// ZDNK=T18GODPa##K28\[0[RDHa<\D3]TE2+c:cAeVI=\>TQ/6X1eZOU[#/@cE;MM
// 3_CAK@2N2IKE(8;S&eS4g<H7dGX1,9;0f.EG70(SVa3baIER8acK,^5[=b&I;2YU
// O=U:M0#JP)3D13H97ZU^L).+N>-U\KO3QB#>]Z3FEWI/N[D.]g3?[-6LYS-9(EET
// 4:fTfKF2_[6]C[)?d]6V.^MT@<A5;.a(KVD]+Kg0T#=aaF5-.+-_-Q_.L_T2[W:=
// ,U,V_-4+<@LTF5<\Q71UQc^9V&gOWY5->^.<#7fQ@CG]G;YWE+PD-[);^PH@ge5g
// T&U-LGMMF?,WOMVb06+&O+#SVU\+3e9O<FLRV4XB@fAeU@QL3,7J+@@RX&N[F6eN
// gV3I2@T53HF0.CX>=ga3BC>H=f\4W0YE]b2E;6(/K8NUG-]93YFe(,Y>T\BdJ?Za
// #-6?&fEB]bMeC-/cCJ#dL/=Gc)SH:/A2\3QIec#@_ga]fN?F#1719<^2[-OB98YL
// Cb>#+>/Z&6.8?A6ZR\Lg\cfZ=,NY1ONda9:8+7dT)f2QWRg<]]&&TLUV@9][^Leb
// /\NQ2/R8YK[A)R.8c-31@_@S:f7J4L02?0CSERSU_dH9@[+,388Mc.HXOJZ+57+)
// gROabSbAYU;3Wf92#:bI]+WTPU&GWCY4Q)OOMDCGL5:AI<PdNR&E3590;Z2?I0GX
// )_6^>F:-VM,6-YFW-#J:5:P@SN:QeQCR-CM+)D7>QT;7V37HWRZ;+TG/SFALfa[e
// MG?J+Oab/Q>&.91bR.-=9;fceOa.=]U3?VggDHI+c44R].(PIbI<BS()M(Eg>6QM
// c5SK2c9^<9G:2LOcUH4JVe9b]#?5PN(#<9>3dBE>52LFCWV3B)Q&fCR^PALV0D[F
// ZZcTAM+<.BbI7K4L7V++:YGQ8b@8E2MEZ1#g]3d2QLX3](#_e3R4X8)XaD0;SYM^
// Z?&IP1aNd.4b;Y(0+T29.NO0)<S:6#fZQ6f3LMV)7#;g>J]14WG:T^;N.0Z5/73B
// PH7</_[B;W\Z5.^L@CaIa2[S<STcCAVKAD7</N7;b1V1SAIIL^P(0aI^<.eF]UJ8
// (<fFK/2<1#W=@=AOOce6@?M:C(<)^CN1@@aa4Y)5?\,)P@JB6A;+6add2RIAgc\T
// F4OGAUf?;:FS1U125&LUYDLMKF33G-O7-YV?aA[eL##K)DG8)6S2_Y/LC>ON?aJH
// H(:d&g1ad5aUHgL+@N>F^X([e(Zd9&&^b&e(/IXYVV<VX8_@]-XJaR[OT8gOWIAE
// SGFg]f1HY\3[.MZYPHCg&6Zc7M#ZWP\]GPO<<QMdL(]&Kb3b&0WFSdLOI#0J7IGQ
// I0A]MV=gF^A0WdS]QPYFcGJCZJIV7SU5eK+?Y4IW?Q\c<0&EZbM1Nd7E/d+ON79R
// CW(2,cVZf4?1G[8>b;eK20KbS3=QD,-VIc/YW?Z@0430^V@^UQ2QX&YRU<G)?LKG
// Y)X<WH6Q@E_I\^LJ[:1@2=.\5g)<4@ADM+1)F)Z7D#6.8M5E#GVgf1Q03F+Cc\[D
// /b3\Uf.:\b4N:#d3J9ZJX6dF,J#e(c.C;,;G6VBHJB8c#\gKB?4=J8CSNGERD0Fd
// c6)I_A\9LbOf4cQ5#RfUg&K:Rb?3S(T[c]_A#+\Xeg5Q6I/ZC=gP091g5<JgQ#/^
// GRA9d>M<^<gY]f/+,=HFf13+4;Ha\0Dc#RgT6f4>a]aa_=b@P@(W=5#]B]dD?a&S
// ME-1M;23N,Z@H<.E+2d>TY;Q7bR\&7gecaZUE+;Na701H/B5.FdAGc0V?.2]#CC.
// EG6RG]C8H).UVeD=#VKUAVM5&RY06[ASMKB:f&@ZdcgIBC[:2J\ZO:.NLWX2ZS38
// @A0cb,VKdBaOPdcP[2_(?/H)V,[YDV_d[;Ad&_@GV(#gP.D#5=D,^(D<7eP[@<7K
// C/=g_-BJ-PQ_Q]bY9W)52Y_D4&&a)>?BJ.HUCU(P7CIW,QM2TBG^/^];LT8_L[cB
// Sb_UW_+D>XU.P(d44GT24D_U]EP6UL^](A6;QW1VIWO(M3@BZY71aGfFd(XZfQ2V
// ]O]c&/49YA,1YbFF[S7TIF:AT]L.?PVI?ERNGa,P#@^\LCW.Z8TUMYXa0J[2)3JZ
// :^TM)V2Eb+_NY27/_QMTb2C4ZFEdbAACRWW3#:W)QYDM>#W@U2QN/=gC#_F)a0U5
// W.<P.XG&3_>NA.2c)A_N4.)dQDZ7D?1E3:U.+;eOGP03eIUP,.\Jc1D#\P5d=Ta]
// ]24/V023O&O;M4-dJf6>&UY=:M4d_EcE-TTU7d0[>=&EAM899X+@BY#;Q,^KC3)9
// D7BOOIfR)BH0_?eQF)PY0fgKBUP>YQH[\-,a6T8NIZ+0Q8.1Rc_<dZ>ZP8X1F5ZL
// SS:HVFf4>4ZTg#9[M^WfP^FR@=>&4QJUHE&N3139g2;?-dSNPOFA8KQX+37AJZS^
// [LT#3E:CfV8E:TUO.-;NRVLGg3Y-7#TK&aJH6aa)TG3K5ZDMD3c2I4\QA#T#gO2b
// =O/RgF05AJII;#U,>b.NO]&.0#V^XKdc@[.?VA^f=QV6,S[D.DBZO-D,M+H5f?Wg
// G@QXcE-@,76/L/L2[K\KLX-H1e)_L+GNYT_BB<7LEZg>B0]+0&E&)FdP&YMeX@ZS
// <LKb1Eb3T1_;Q6bKeXV0Hf]57;3-7[(1]<X[9cCd&8c1A8CZc)>O3ZMPL]3P3ZZJ
// MOdU.M>e^8YbeIdW-\7&U(I=GW3:NGA>\Cc?#EB@5]+7BE+@@=YF25L7\HWE-5&\
// P9(8ZD^/P#6Hg<Q7/#L8<<40I4fI>ba#fGBVUfT@4b/d@U\3)J,(dS3H+?D@:#ZY
// dWV=V4a57K1EP5)^[V<5Q_UJ=>:/aSC/YYQe^deYTFa<,(R>1E3>1DY@A//<a@FR
// 6TB@EB>0cX1>d3(]&\MO3Hc>ZPg3]dQC#b#TZA:V@f-2g\K3dFNNF6JBUCB);R-X
// DM+<-/QMRL_@eGd_JK+(GeObCDUCf)f-T(,6D>W#>,73;;c\?J8Ue(??d^c\&dHF
// &PDf(&6XG#-,)[Q+@cc5Z>Ud3d,Q:A8:9FA,/H@/PE+UBS;I4e__8c\RL5F2EIQM
// abY>YUEWVZ]BH,7J)5b>g391VbG0.DX.^H)6OZW9D]Q>WA0Cgf^fHfKRTg[A22X)
// c/GD&VN<#(YV?BbP/ZRB^I01NJT<9-]f9AFdSbSeGaY<RP\I<BMDUHRL5Bd)Wd45
// ;;4g)RB8UBPN&?I(D7KI>c?4.^9+HG=A&#bc:X9SSCT1EJfeg^ff:E\QKW@<0OH+
// [4&<8Cc_T@WZBWEdPOM]JKS(Gg\ZU25A);<EE73b,>,CHe9[95VC[3NGN@JW-LH2
// 0EdZ^H686.5=#+]@SaCTMUIENNS.g995JaI?D0]#NU2Z8,@;C]0bT)^5V/VX)FB=
// VBY?cJ#ZVW;G^;:7WP17S,LN--)MO<,JeL.]:_;W_><[7g:eYg[5..G<HD5Bc&Ue
// AK_;2K:LVMRW>B/5B]Q4bUA/XMD-C-/dPdD(gC^<^d81G1[OVDF3>6B3EU&MJ=4^
// LR/PK7T1=aKRTa].<MHAPRW15]W5(8X+;DSS>ecbT30_H@<M:?#e+N\fK91Q2)FT
// TeNQRV4Bg6E,8\fc50M#^fEKO(;?<N+bVe&:DG@&W;<6:GN.QN[c9]a@,,<XTZRN
// 7B\6IU,428a1;KCZ[:6b,3N7TQ7Sf-A7\)D+I>Q;M^cVHKS(_(fJJb#7N2H?gc>>
// 4?P;G]X-1Y3WF^7afFKMYeQ_+&aHS,eXXE]0gN:_WY8JTbbgDAVgG9Q:9.C07<G@
// )SCDa,Dc@F9ND[LW/Y)(V<RgD^2eP8W=XL<d,/2:fV8<@,>4e>^G<c7@3/S.W\D5
// 7ENK&44)6ZTc)R6?5OH<]2_OJ8F2;FU0YF@^00,;7ZT)5/Qd>g.7GM,5gI;7VDfJ
// 5@_,d?EX88B4g;G?>?2ICP7We:A-BWUMKNb@_-6e&TQ<Oe<#PdG^LNQ[WF?8EGA#
// 6(HEP?LV<G>J.-A.4I9gFD:?8cQDR=&U]&N.R5Y(L&(WdHcHV7/PW:]a_#QeL015
// JWS1\T^]U-Pa;]3/25&AdQa/ZBE4LT.JG-G2-c2NbgQHI>@W[_cW_A[+5F@,;dOR
// :J&TJRE9DAFR8920b;W?I17N+<gRReIKA(IOXfcX<?E2CH[fW\Q<V:7HSX9N&UGc
// J[>6TcM:A?,>:XRHc?LH@73,OSVM#:SLE\7=4RLTe?YR^4A(9:186VODUR,TZ#WU
// ]3V@ABUKdH:gT&>]gMW#AC_aCRRc&XLJd7KNfa8MJR@FD&Q1a9&<#4e-[+e6\KeX
// RD_[#>WgPaG4K=YI^(+1b\(\L+OH^#M.=XDS0UgLeg8(UU2J>#URPg1S]#/e41VQ
// .\,+4(4T105U3a+MMbA_SKCc1=(/e_-510_LO(d-E.@OE.SH-#GO)E#eVUJ5aXA]
// CYYOMK@_0YGACRPJDAcMB0<HZ9UV]6(+25Z/P+A&9<()1+7.D;de7Z1MU_b#<aG\
// @DAYV>J2[..)=#,T[TA7?_dAA-QY(J41ae[Dd]Le<QO&;30=BI@[?+c(R2?[516Y
// 7D1A,5U0KK&b&@@,WE(VBR:MHL&AY.),@,EO5BH3SWcF92cLcCTU=,@7)[JV;/M]
// <Zf1BFBHRM2/a4=PJKEQg,2422(<]R4UD?-JAE)Y.YQA.eK.L80bge<;f/a5XV_(
// 34S)eb=WgAWZB:5<N+YHKPf/gfWfcLX>cce]e3_AIO2&DbER/E/K9NBd^LDa3TQS
// 5f0#XF-e9,dLD\9e83/eW]--H=CJ[X;89Qc0IHFGcSX3:R_EPgCA1d3[VX6/7I11
// 7ZM)f@&M1CgW0>Y@P8)g^ecOIPG<@N5<a4X[O<P93G>.1Md:+e=,A&YUP_RCE8T4
// <d3;e@PCT<6S1SB9D#T>G@M1dB_2@,[>@(dW&fBI938&[;B<Ge@W+WIEef(04RR2
// FKG>008\?9=PcPY9+-0&Z-V8,a>X6B)]6IH7>V.&J;9E2d\R(XP)@7^<&3(0FEDZ
// c)Yg9+(/Sf-/^=B\J=LFF,<6GMY8W)e=54e\V,-L1eQe&O30_IJ@D4VYWHbHWZZ#
// WfOM+ZBI4XZb(Z2EbR97T5d->^,=C<\gX:-T&CF-;2TA;)RV]BN<S:VI8UO5&f&d
// ,EeWES]FGa:32=#<.;85(b[7b<a;b;;SCG1M.Y(c__8I/XB6ZP?\X_4Q2PEZ7/Z1
// \2_)35.MdL@McZ]JHD6^+Q9B,#G7NeIV@1eJHNAPdd54Y0HHZK^;9D888GX=R/A4
// 1WaJKUH,@fVbb.J\[L[gX.)RaCKRJ5,9,S^=;LZU)RV_a]J^<\&4\:gEJ4c&-#[4
// OHL<@@<NGEP=TG1ZSX[I;@=EOW427Q[;,@E@6RS<LDbbRb.^/5&I+03T1V,>[6FC
// _]K.[N0VK10<WOGV5I:gFZa:+SHG^ID:28&G/ecN4<U6J,6G82+2MQF&@TS[TP3]
// +,_Ab8&?/ff^Q1K>EcOVO.QS0QW;PTW.1^;R0LS-FS58S56;2S+79AP#I\)7@4_E
// g<I)I)23Mf,caTBc(X5FHPVT-1A=11(/6d=.c_P)M@Q/0B0bXYWg4SL9=2E2,(Wc
// \@&JS)&Xg9QDB54_A8Jc9(;[50NIRQMVIN)UCV#]Sb?>9>G.aIK(=#,BU=IQ00dP
// F<&7#L-==Q.<N]eT,XZ&=6J7DL(C0#LSJ2W(;GTRfa2964cIgX1W=49]a+gFT5K8
// Z,93>WX>Te;(1[gYc+.Wc0f78QTb3-2ZcEH/:J=&A(7=4X)\G^bU.,-ZOVYI6_\L
// e7,GY-GD88J5K<F;B>(ZHPSTQ4VP\cEKfW?X4^N3?4+FI_Dc?dO?KUV:KdT[2[TH
// 9&7ON#;ZNfJF4F]Y&X,e[b6+7aM/WXLOZOQZ85H32IQD^3#:#c1[d79CbYVAR/X)
// ZbA:)I9[RQJO6YP+)P6LUGQEBZAV[20_L.eZX_B<,GN]UcOCN\Vf42]/ag.4Z6WK
// f+SHGVCM[Q>+VfE9SF]g<CU/\YJP,R])H?.H3+<69032ReQZ;UG\N+11fTdB>H\+
// b7b=\@@36UUFQDET7^O5PBC?#\:E0/=V&fA))5Z[dZ9VXBaQ7TSeE?UD)@S^#+NO
// :\7E&d9;;0UCK-7fHUMVS5b;TG=4d#W>9<9@fD71I\4;TG&e5H3d,(aU>[AJO6KY
// J_I/R7:bR3VMDHBAREPc=IDBA0X5\##=#I.)<Q#/YEIgE\ZcH2d77fJ-;RXB82=+
// J89?65E9F(IS2KVM].HT27II&9&M&/2;;a<2@gbed_7510/8]@_Q5C<=\O3D/A12
// @S._@3+V:M\,1P)A2<X@\27VR5MS>0=9]Vd\ceKL>0#J0SCS2E2c/RO:b?[ZD,Z<
// e84c(U1QfCPHB#=>\eVEO7<daFV\J76GE9>BM@2e;UaCO+5&Ke3dZVC]DdbK800\
// 0=X7J;V<.8KUUV]^D@1d[U#\dDN#/^/&XcT9R^^Q(#)TYLYQJ63U\&eL@W3;Df>U
// 50M[7(_IcVMJDB(c]KC;58gVXQ2Z-[)^T:EWF7(bK-Z82//EIB2FMfPXU</6c5V+
// dAMRZ<Pcc+9-))YO60>;Z6UPV2PRSfFW@_2]69Kf,a.L._HJ>cc;aZZ?[G-MVPa+
// 6KBI^/YA6B5KL6DD-OdR9Ce(.B>-88e1A[AHW)\1HJW-0B&f@\-KMY[d;5_5GcfD
// 6=@+TROKG,LO&bM[24D=._a.;DA9I1d.5fdG2WEF,]4.bc5>YFN^]MH:(f?0ED)F
// &eZ&>QB:P&PcYdb9ONW8Sa:,:..EO4JUKW6KMA=f+cL;&)<MDF@RFYV?BO?(N0Z2
// bD5b^:0\Ec_2HfRFC<N8R5H(O^C\gDH2>CI\9VQaZ:2.aC53+P5/UC#WZ/1TKgN<
// M/TLF=OGQc0G7ac<We4>JEfd5gd,F0?gJeVZ43,a,VfFD\.^=H-5,gSc.4eD0-c@
// C77b)FCR\c<DUCS[&J<g+.JE\K48;G[d1^9[1.be2a9,HW1U4KW4SfPAa6-P(d?,
// JBW#fd24Qe2RK1_/#?N1,))6>()E730I(-,H8H/ZZ^J-c@?XJ?DdS14X5P(=d9H=
// BbG:.ac&8gYI\Y@6D3M@MVO/b_LL#ER9Q32UU[_0+G@\^,RNfA;@S<1:U)H_#K7e
// R1\bfU6Z4.)_-g-Z_=#.KQ9^VT+(>241X@GRM2OI9U\]>I,E0XA#Z&IZ7_+aSZcO
// KJW,K-Y0f\F\7aW]B=B8^7F^E]/O+VH<5\Z>d9eFW;BNJ_<>&gaC];,<F^L1Ra&+
// Red\@RCaT<2X)=TaHF[,e03,UW3R;fJ-@b/<V_PaKeIb;.GEF?XVBgF<b>P=<C#O
// ()K(P#aP^XQ7McE<V9@cN0RT5CPWD]XJR-.d7Y>09XIfZ<4UDC80H/GG-/1QGK\]
// R^GR.H9>^9=C69<[PcV927H#dT@FMBeT34,(VXFN2NZ<<<+YCMR1b0e>A<\I]JK]
// >FdeM0N\1_,?e:gTN3g&<gg(2\A&KPNAZ7KER.?C8W4?De.BO(]?BHX7KTEJDQf-
// <<MY?-L(^A1HF14Q8U;QXd1EJNNRO;SXST@V@9?AS6Pf/Mc)XZGD&[3#<WZEWF@/
// S.CUR?4R\La0T?/C4g(#/NZ_geUagBG-UDSP16WL.5__/e3T]Y4F-d]-G@GLEFKD
// PU/QfVOcgNWgK:f@KU?HgN7dXbQXeBaR<55SH]UVKI+>@fR6DY[H:dB]\VX(P-],
// V+FHJIf,Hd-OH;bA#@F0@[b5gW8V1&cM:d_5HN(CQ/.YO_dQ.9),GWI5&9aB.\D=
// IeYO[+3E4bH^D)-XA^V?+@MHS/93#=.5ObB\+-\0dNOGfLf6C&E1&-WdI3dSLO0D
// 0]Q#KCZ#<,>acN+>A=bF_;\LY7PacY[bK&:34N^[R6g1_F>JU[Mad<OL4UIRM&HR
// Bc-O)VLD[-E]J3FP/X\PgY_F.(2<PPR[aQ)J)?a-821A.2,Qb;&+56>3#<47(2<U
// CE_UBOf@=9C]=fR4?AfPc_\JgJJ3fDb#_UH622RJLQ3:1#64MF5&FZFeDWZ1OHf8
// Y[V<e-9=AGdb.+A)#a7:>^+1dXR9e[RF<0(E,58J2M[<>;(f23@5E9TF_TRK(;[7
// 5\E5#a)Q<Pf=H2M.RQC2P&8NNf9G,@;(^9]CFS0-DXfKEU6Z^V<g__)\bN<gEFX;
// 0\@:JY9AMVMI\5@^?9QgPC7GM<aEQHcYbY.,XHDU76J2L/Ma2g8)b__3EOag3S[_
// _D-92&Z@a-7aP9\7a.F/L=L3,-ML?J.WV6bg&gZQC>:f_K?[33I<[96P<b<O?[14
// 3/KJK6AN:&J-<PDRWAJ6,edW[MH\:28ELSNE>_?GFXU)2J2bDXc\/-V=IAF-.II6
// \D44(&,UNK(bd4[N?BVef2]dLR\V_O&dU[.2:GKA&35.)SD0<@A(H+I>UV5>/W@#
// F;e)Z8FX2P@OS+9Q;O>Y52\U3&D&[LN0IAdf+OK@-S60IQO-L[_OC[WNQZ(V65JD
// =QDC<ebQ[/W9dPgDfE71d517(:e#dS<-KK=09#IISB-G^[(+2fWdU#:dL,E(<-&e
// R#f;b-a-=M0VY724OQZ/,4S/M>5V8;OJef0#g,5A+=@D(Yf=_@/TFY[DB^G)A8\,
// &W6XbXV#YaT,E37AQV.EdWA4J.U3Z5^:=E3&F4GW\4XaYVPb+=:aeYD((-gO#3Y9
// G4?GKGgO?MP_FcTU#SVY]_4PH@KDQT7YONZ6\aQ)2HVK1/?.;RaI_g7cL<dHE<QG
// 1SZ]gc4B#IALfdBD6<OL(:eROPcJZ5Q_QN/a^YPW]Q?P@.9KT,fG0B23d)2OY<Xc
// 9V?I?\//4G^=da1/6&VZ4;Nb:&>4(C<@2UK[C;OR52d6D6_8>V(S6QQ25@[8R]c)
// ;,7>BJ()LM^5E[cK5UTb+;eL=A6@dL+3F9cJOKPS<T7dN7N0G>]MJ@/(;MJ9eTbe
// #]@W201f>.4cHBfgPCa,PZ<AR[)KePZ9Z,/aZ]OU6P0EHQ9^/3eUaB5gGVP1VMN/
// (B=geY,S1>70B..?RZ9&YY8g=V^g&W[2X5RFX1?f^:2c0e/L<VVJ,@XLM\),I7#c
// #g1QS^,FD)V/(Y=,MGf>f_&<KE5dXO,<dJg53J6.OTJ#fMF^VD(I=gAJWP&FL=/2
// 0\[?g<fD\ORG[R0g3XUO4af5:cd,0Me]]W]E.9MCg0[:^aI:Fc#&Sa..0Xa@D2]H
// \5(gCH31PNAg4f.aJ5;YBI8?F>eAB?V.U(>:-8c<PWDN+BML;Z0&,?PWMOBW43IX
// N5HP&\.>EQU[J+L/A.LN9C,>TIO)J1N2A(8=N5\d<J+@9?#K;)b?d2/dWX]&cN>1
// 21>d\2Y<OA#BV_.)fgDI0INb7ecYOLT4)X-@RNILC/B&W,]1#F)^F)0bcA_cZZ4Z
// ]1JB6SUXN)WU43M,]H;@E1]_NOX]TUd(M<=2ZWfV3B)^fD\)UW2E@HR\&^2P?K7Q
// \7G&+ZTS[T.(Kd4[<79[A[B)aZ?FGb.\G@UgTd..36JZ[A/U@&N0_>5E)1XJ0K-3
// #L.@V[:;+8<+CHN/caLCGe\ZNCZ916ZV-]<D(_-)<M=])HY_VOEd><4a8M0)dX24
// UE+=XX?TJI>H>XI.gRLUcZ@Ia&LZ7@>MYX2>EFTYOGYCM-5E@(e2c/OH^.ECe+KF
// 4(#I6d=W2O]=@),DLQe.Ea;HdJ8GRYMAKJc#49VNY8,4(JHP4R;?3OCH,IUQKgF&
// T\4e9&LcGHMBZg>_RVfNUTf,X0?gK/(gP.?)#,Y(&N16&Za<7LWdeMcUXb;[9RgM
// AbJ.9[6@N_]a/RC+5]16YBP99SD0P_EG8&.d^U3P:)IBb\@93\57,JLL>KB/P/fQ
// /KIb2,X^g#ffU[#Y(N:=>PAZfH=N)FeWE?.R.Qd?CK.b5L1-VT9cA)N(@R67UI.8
// e#Z7I2H)=bd#W9(GYBB6C,.NOB&eQ1RE2R[<Id88UD\0V>@f^KAG:1U_S)X77MdH
// RK.<;4G?_I#K8AQ=XMTGdE^V8X+XPE,?O]?GL>>,a_92[ORcQR.BFK>.Ta:/X-]/
// \G>B[BU+Wa9]F:XX96P9,M6(@VJC0#V(VG&R[CB-fReA]LLN#,6c+UV\,,[T6)7X
// M[CGgfSa6QVEL@J2Q)/K>5]+#@.N/aFCR6CQDfO&9C3KAICaPF0BLK)?=C;V>HSH
// @AZMJL),,/H,>,2bOOb&S<aC66L-578;FYFK]F?R4/aAR/X#2C3bHeK[X3SP2^b[
// _[PPb>TE51cT:\C;?Rb/3O170a0,CUe6Ye+d:&Mc#b<YK-27#9)N;a5]]<D-87H:
// SaEU4M:.K19TCJJ1a;Q_;b+3V1:6bb^dbXLU_Ma^WOFe,Q@0R9fF6aU1O^H.b.28
// 3<-T-RH8XbA2faJGI)02/3Q922JQA?8;g9)N\AF=1]_KcgDQ:;/Z.GSH@O@Z.1ON
// :U5&/+\3:9,I<8+O6]W7[\X.Ee6#E03fEJY^Yc=KWb4I;]d8_K@L2Mf8ROIM2dY7
// LIeSL_YO8LAY]LMS##KN(,L@QXC:/B.&:[^g6TfA+T4>V#/K>Ga#b20W,2^eN0cE
// /0C=f9DYW,1?0?Va&+)[6GgJ6K6@MfeG.GZOd\-Oa/-gF1aDH:XXG?:W+eIO&(=P
// =HFZ5^(TT)4C,FU@K93aU8)61gCACT7,]=3UIQ1aKZ+:QV:b5//@d@UVQPQ\Y7]K
// d(74GEQK/RaU48.^W/>:baB^C-]M/6Y-]E6&^I]5,fF(Y0A,eCRF^AP>1:,b\T8K
// 8LV]BH5OMVYga5L.CIWA@g8B6..PM@-K.;^LK+>J_.f&[I.dMUM:#ZDN;Y0a?cc6
// ];@0GKZJ:b#WRHE>P=):B<10:3?2R\:fM(U8L1:8C7G=TKTY#^E8g+Xbdbe70IEg
// ;+H_W-7fa+VMVFM6c:8QU8<15?L0E3QF\=G7WU&(D(KXUE]E>VgYXV_/gG5KG.+R
// _VFI#82=MU<8b/d@?55G<gbbPKNOVWCBgMc91D)KUd-6;9EG4N:X)bK_R/06#Ig0
// e8W41:Z#Jf]<bJ@/(5U+6;0?8:,?ABBbAS&,bCaS9\03EW[1KR.>@+/KL:IEX>HE
// /D/A-P0T+ESXYW6=D-Ve(MT=.(&ZG(LR]]5N;acGS\;f/:&^AV;gFC=7=[B_YL#Y
// :3gFU(@MKf0\E2&F6g6eP]S6ARBVQXHKAFR)8?K68ED4<23R]6]OJLV+K<J>;?6C
// #PFJ8<V_+.6BO7RcAXKd.6KKCF46N3VTfCB@46ZSZ=^(_;Y==[/Pa70eV72]e><X
// aPBN.K^fTUJM#&&IfI-+9UFO;T6aB)HYW,N5_7T#GX=>_U_/5C\?ALSX:A<&GU<g
// A;B>FX#@K9WV/NXeHN[dEe.4>2<VX_eAe-ER,/(U1G-c2L6^Z9>DF8Zd4fa<,_=S
// .#.U./Y4.U>/EHB,CM3\]X_77F3_2#.@QQ+ASQQD[]U+?Y@##K)2O>2Xf]S)P2\:
// K^@T/eMffC99=B-=<BaN)C(5+ad7P<BHDcfX@I#@ba9]<XU/DC#DPe5A:F=WX@WL
// CPDS^A5HdAF<AbJe0=Yd8dA-ID]3e)RE^J\:9aT33_SCUHUFSaC3@RY[-6bTGW(Y
// De_c)W9.dbf+>CF@IMB9OJ5>KZCH;Mfa)KP/>7JUR4+(Y2INR[bG+N8fI-1[a51F
// #=(<M<0+V.XLdYVW^?<?W(9.:;Z);_Cb;R3RH\PP0Q\UYb1P3d[S6C.5S[HI,1eW
// SXKZ^I>=;fX2c(L-d3M\6^S4+6:4NfbS\PX-4ba.CS-C26J:GTT6cE]^3[?g#[NX
// 0&^;W]X>S\;PLP&?MRU<DX^ZT#c,]6:H+U<N\:fOE.TfJ(GB0TR,H2;GWBX.62M>
// @A>V8b]ee(R8X4e((+&2HF\N6g_>^+N\f,;E1\J&W1d[^K>fSHKf4FFE9Va;b,>>
// &.:EKgDZ75MY5H1A;#==f&?=4ZB>Y10WRD[DL]8]Y>/;H@_b<cLG1TD^+gDde4_C
// ,8SJH3g7T;BKTYLR7gV0#WI;PZGF.22Z4-b_?Y41ZZI+U/R.NX&(ZA/d@_8;B]+A
// >.=4CHVG9,VX/0L<HJ1F/(=_;(9YJ;RIL0F?BRJJ@:I57=W[WX,.:RY&M>7Q<\aA
// 3cbTIV^9dEAVQFI3:&F0eYg>@^Tg\]c9fc,P^b)(gM/I>L(-eV<[X1F,HSUgNE(T
// &E<D8]4eLFI,TY1Pb+f8:J=87GE56Ke(^KQ8BD1S8@_6LC.SUZe]YTBaC7O-Z7S1
// PHGB[2Qb8DU)#?We<M)a2/Zb?AIW))8D36+C-]H-RD?0^\^MgdIS,,,+ZaA,52_7
// D4C_\6C)N:LDNLT:72BO_Z3aH1L@cV<W_88aA=>L]&#N3V?;:-FfUK_aPcN2G2P1
// )X)EeWX(RAg)^<)[7,cgAD?>\B_Z1:TM)Jf[E]M&g_05G[O[)/Q:^7ZND?&<F:d?
// 6d#XUe7cYV@^=T(>.QdM-].9gDDMRXF&A\FB7cWPN-BfQJ7KI:Bf5TG:DZeJY;W8
// <UVJXD]?79<Va:dXQ1#\X&RNUU,BVP?B0WO.4.PL;cN>KW>c#NeT]Bd4CGNc(F^-
// S6U&9G>,[8MCT+:&RZdO<P0>^b[&:Sf12?O4WO-4=X\=,HRb^?MgY]J@^];:L6c&
// Mb99cN0W_L7e_)G2Y]dfe;;]AcdEPC@H(2a-UA]D5d62EWaT2U(/8=,MB#\1X.<J
// 4=CEA6)C([Z/&=N08e8\B/L]VZY11N+P8b:\Ja?W)Sc?+g_F6[?X1&5^J^;Dge2c
// a(;-)Q]MAN9N92NI#NEFbDV\P0UP5M2@S:/)NB=6c6#f9BW)D&W8<-e\&AY,H7V-
// GbTZ91b#3LU0&N-9_Q./DYR9gY<@IE_#-SZA__YWXJada9Lb=5=ZK7PQ\<2g[CZT
// 75MPf9;6EYd5ZA4D:SZ94X0LWbG2ZV?D.8>G+LB;;eOKK\cBGSb3U]AfSMK_3EH_
// Y4ddgCO5SbH);H&EERRa]@:6^-S];8B9IR]-5B=+gf5:faVPP2YO=SR^\MaL-g4H
// O#)S:a4bD&bY?P&e:9cRE9BGRCbQX1.7ED5]SOc]g-0O;SNZ1e5L>)BdVNF.[M&[
// NE\JL[8#8^8MI=Z8g4Y26fFA7S\H\\Y^aa:Vg.fcDg+_0bKER6:b:TEdNM(HXgY^
// 7E&OI;PQSd9(R8T[TCM87WGbG@H\(8ES7BNRX):G>E2aODg6d2Z)ZJdAB4Rb)UV-
// )F,gMRb1(8C;2[;(eF8QG4V?(c:C^:dK#T7,PA#GYBU_edT+56RKZ5eS0.GI6;V+
// \OY/:R,@\]_YdV<:GLR)bE;K3-0)Y#1TBT/Z3+9BV[a4_GXdU4WL0e\J#&4<)N0.
// <f]P^/KD&\6ge2P(1fG^Z,EOX+?GO#T,XEb=7He<4#4U3#F.@7)K;Y)g4c;0VcGF
// 8-8KMf^67/XSb0L>[bYgQ,&;?2GUBde.+)+.?:IBN4ZQ?GZaWeE&NZO<&L)3]>,<
// _3IOF+2ScZe8=S4/g,8-(AHIN-3B4)dO3\9K8Z_/J=9M-=d#b9E;I[C4P=;WK[eB
// Ba0WGB[^1N2O@R=N6:-BR_B\Q0K:CWD_<XM/:Jaa8d3X/fIL&TcN68Y>TS:eA-ZJ
// USGe0H4E@(GV?LB-L-+127gH75Fa04^B[Ecf=@P]W(KNBI)73ILAPWbL6=W2g4@@
// ?2cOMWL.8gX0;b^)3;J6]=F^&>6AK#CCP6-MF8I>?13DU<P<Z>#,dafNDI&g51V]
// :I)HIDF#7Aa3.cL-7:a8K;D2@OA,]7CF\1B[0._A[>_/FL,+g;5D<7[1J#EIG,?9
// 2A@5Y\Z<Q^7I;Q([UH#98#J8:5FGSG(W[@R#+4P/TXH@b10a]A+Y9W,2+KdMF::K
// =[96\#NbJ8X/7<g<WZMB)cL3#QU^5BK6?9Q1-G>,D]Bf>HcM>Z#J@0<DK0)#<Y_D
// EV;2f5eOaF/PVVJI@W-CN3d12PV?:F.(e?\_GFg<?)bWST<5)B>>^RD1b[c_+-Ye
// &8/7Y#+#T:)&9U.FVBY]5@^[##,4+G8U0/2P9J,K[1CaU)EcJUTYbfQQ\FD+I:8B
// K<9IHc5bOQ2>(47NXNZc^5-7T>dVHK,#IH)\R5-[;8@)WR.KdS.T82)N(+0PNM<+
// 2<J?>cY_I?5d:,O]<FHSKW_]gU)(gK(<5G<(3X0D(gR)/5gZg3@f7A94[CJP_2]g
// \1FFJ_)#5HdE_OFCJ?==:Qg^[&4EQbV_@FM(SPRDgFbZ94eI8]R.OB&AaRR89^>S
// (e+MLKU&S,T--#P0.PN_\<)(M&8AD@8\-D4)d:;^4:@T)F5cP&]VYS@O/WZ_fS#N
// 6X[@=/c6Y/fI_QU,>^NGFFW9&&BECLS))[[2G,G-OgFW2[4B853T4Z+LV,P?I&B3
// 8b?UZ8^gXLA?JEf6LK6ZR7\:AI-Z]W:Y9c-^KZHVWNC:PN_d5>a66g>]G-\[e>.8
// 5E+aZ\TIT:(D#K\/D&K^Y7D-@a;?.11,780/;+0..9HZ=QJ0Z/#]FF&\K[@>d=M1
// GA7)(<H27YMIS?a-&>FM9cdBdIWWg_^[eK1Y0AEI<.ffWOC;&c4KZE]1?YD4XF9>
// >_U=dK,)/TCU0[NNFg09G_e\e5cQ)Dc-&KgVWcXN\36.OI6SWI9Z[N2W\V8O-cKT
// a3>=@9f)IHNAUFc<7]b92P(5A9VL[G:X>eGV);I=]R:/+)UXIOA21OD2;8[_3e2S
// 7aA61\Z]1)Nc[1OSZ2\Z@eFA>cdN_W0YJf(&f=W9W-(L,-]c+P]NIf&N]6UH@US1
// 2BL@Oe5/QH9<L>Jd]>e6.R#]C_>;OgR#IDW?dQ#+/S]IU#T4,.QKN,.V@,)d3#/:
// LgY@?C12\D2AFOA>cP3@6-HGbYQ:,O121-7&P&>Y/5N_bf?JXK(XZg:CbgQc=+?5
// B<E45T0PW4dMg2<2(9.27F-c7>ALWc]c6^?9Lf_2cNNA\CaF&T8HUHaG^VJ;/,/Y
// 2b#/91[VCY43gH6UX#cWffc,OgcO0/6[f@:3>\_6S6>X@\^g=EOK2-P.dgCH8D7(
// 9b<ZDQSM>;277aBJQ>fP?LY?_YT>L)N<[cP>[bW9>OK@WM7LW._]6-G2N<FeQ>2K
// C.ZJW\a]8VHPXMge9=F=O30gT2H<(e?f=5;P\?HNW[?-Pd.K#f-4\ag9+#P;e/4<
// Cg@#N?Z@IcB:P5)d6_BV2g@7&IKYdbM6g+&R@CY\C@[+:LE9V(/gIPI5Z]=B>(Y=
// g1TV7LH9>\GV:AIB8Yc\Y=NDB?RTaUW_(PQKdV=a3[V6?2:\bE(19Tc@Fe#F7]:Y
// AL(Z:W#Ud651:#[e(aK3R(SDeaS#/O@6__)O>Y8-AQVe-:&DGXJ+:O2<VFg//B&8
// @(N4WAT,,VWFQ3f93.3W38Sf,+e9-aOdC;F70J=DT,HCgaD0F&dFJ[0O@5N5#WPU
// G4QW#TKMNE?WfD.OF6QH1C3_9db<&Y>;?HT:d3/FD.6;FLV90XWCI1/P+7IX(d#7
// N0/N+(QENSYQTWDDcZVD8_G\?cLE>f/8(T6OXFeK./#N:<P5JaVFa@F&;68H/EL)
// fa=#_ZHbNGD8RQE/gb58aO1>R73C<1eNR)5g/X<Q1JW;TE5(:Ng)/IXQaK]=SFO4
// C-a;0O45,g1[K:71WBC=KOYAG0L(\)#QK)=R-W+/C19.OUf+a1LVN1^X6/P4]Oe=
// M12b3U\,KUD^3KbLE#LX(E:ZTF8FV>Z/bKJ+cFe62/&6SU5U?1gf4RZ8K)_M.88Y
// BM=W_dX_TM]fB]g.O]-2<:0&Y2_7I#7P:^4eaA,UeF8;)IAX;HG0#<&JV=Yg^0X,
// GR-/Jb+H&7<?LZd#[KL@eY2R?6QY8O:LD/1H_\>L8c=>QG915@?fDa\4Ta[Z;F03
// 1\H?8YE0HZUfL[#6@G<cDTP;1K)8fL=Pf?@<R6/_Q@bI.@:7#<faZM_B9_<[;M#I
// Be39f3_G4M/6(Y2<&\8>_RNGc5H\2g1:]D)#ZCSPAMd7WII+T#9EHO)W[:RMB1RU
// 7)FB#FW\(cJ(O:UHGD)V4J:R=Z,G&=,/_TEeJU=9Pc;O+N?Fdb#FD.>d=d6b,-:(
// WLT0O\1Ze48S0J.<<_S8)P^EBDY[5<#/-EOX3<9Q=d#UFP/YZS@2M58_5U?5RAMT
// <cAO#I)^W>^(@2e6([dTOY5YS^fd?WdR8IeZP;WC7Uc:5e7(fM_RLf7Y+II>#4/2
// ]X:PV(=_)DT]70227/.Y8:C]2;/MZTO-M?O83NW:D\ddNgdS__,62Y=X.RBbK?0V
// b-GQU:NPM2W3/71]>BM@/K0UZA;=1O+[MMQX?_5Q?<^]F6g8Mc_gQ\SBa:<N=?fC
// Nf2GGN7O&P]8MAE.PAYHL1LAJbHa#0X8\.aTc)SK#N-3R1US7_d9Y#Vf:]QL.>::
// .X/Gg4Q.a4_AT\,7YXYD\X,PIJUZ\+BgEB)@C.4@07GK+fb]/R6VP\SCV&\gKJW?
// e2I&G8Oc8+LL\2^7U;]N5AGFUE8X+#60RE3T[#UgIAPW3LJ.LR@U(9C?&S/AN736
// /-F[Xe[G,KF]+\F7cSc]8VW)-=1VB//VZV,0WFLNRD4CK6>/+KJMHa4fRUd90U4b
// XbH\Q(_(UOM=c+2,W:F]eCV?C.\;fL>g77JU9CZ;g])\7eTbE0);XPaFXQ]Z[XKg
// NAENH/A)PM>R<1Z5X0\M._0^3KDK.PV;75.6(?]#[)])?C4<XcTbIX&3Xd_XAQ9Y
// 8[0X(=6cfNX=<e:W+Q7\N05SeUA.HS:SfP+9ab.406U[OHOd20K-1b^e0^Md+=0,
// W)0b1)32Y\)cE_K]K6=3->;;.Z?,^_[D@fF9_d_1E.UT,3.P>;g2a.2HSH[>[2CZ
// I0Sc,Fb2UG=\LD2SeCeE1e2PJaSX90F1X7S/7<,RK?Mg_W8\-&,W#6+YL,IKT.C0
// X3RI7_T28b5Q[.)fe-LD9J/8VE6X5J5CD<BPa[9Ya5;0cSg:D<^W=P0H1<DH;HC:
// DOC6JJT&&F5&BQa4T.5[fPgK-(,A+JK_4<Z#=J@HHJe_+O&BIOTE;[5O\H#de,&b
// ^8B_#\1aS)<7Q23:>^:1A:83d<]EfZNDB,ZJLg_SKM:V193bABBSB^[SVb0?ZK0N
// _,?8AD:++O3?KX6g8P/H@?-Q,AS;SZ;bW.?^DR-OdUV:LIEI[R6PaQ3]^2(&\A^-
// I^MUS4TbZZE6Y0S\<=P_M<ece&dEaRJJ89dc[B\QU:WIS2a>Z&X:aLR+6#2X;JQ1
// <V+TagC&TGB&_cgd:?,7?5A2Gc-JM7;Hd9]2?#UD]<TE4U-cgDW4E&5(a9WIfS\U
// dd5W=C08N)DC7[6+];UMdb3^\#Q@2@RCZ<LIfe:E.0.S/Ef(O?]KC:FMSF3:J3??
// ,TKbX:)G_&[)STIH^=L.6.a&PZ&_IQHQD0NC(/cH,0RbPE.8NTII?b)\]YXTf2:F
// J.(B=\TgJJKR5ZcfT:f?O)=C3eBKT_f,.8;627\c)Y,IPJGZ@-<gYc[?)8/c@JXg
// CbgBP\>BX7MHPR?/-+7VO_-2WNXNQbZfF2V_5GL[Q:Mcf.aWXNAP&R4JM6/0J0.6
// CN?Kd#[dN7&f1):@QRB.e_C]\HEE9+3E)NBY<79BL(P-M9ETbW&Zc?0B_=/8&OT[
// O]+V;#Ge]HZ37EMY[\(G7V#-]eP3)4N7c-b+1bSHZ,3QD<f69ffX_@aEgb#<L:Z/
// T1/QN=#GP7NNFIfd37W]O0TVF1P6;[)L&=P,eG;aB?:C#)+SA0_Q.6782?9HKA5b
// YOF;&I<c<]E4<(bbY-V7[,LB),4&FAE)e>M[g/,;?ZO,EJU5.I3OF9cV?/L+)?0P
// I>9T8PSBb\-?YG(J]DFWL+0<bTPA4K=bAMG5JYP<77^W6^-5./YDZB<9T8,>F0H^
// X<31&E<-^)L[JLKL_065D9/7L6<I0+E<Eb[N7Dg55)WdZ60G[eGWO(Za8G^0XOcV
// 86(7MJWeLA^]2g6_UED.f38EX]d]4B35T=1aOLg1a&:WY0WP;&ELOU53Na&fB\d3
// ?PI^^,W[PWOE+2<:N2VH0FAO&Z(=/:bR7e76T63]ec4S)(N63:]U2ASH=RbO>M-1
// 7)dA+T;.gF62dg#S@Gc5?AA.\e5Y<YH,G]Gg=V4VF=4(<H>agdMDK8M0^..;N8W5
// VbZ:]C/De9:,d]DYP]AgAJO&5<<d,[T-N?8LY86+e[_YX]XZ35VP;-^R]Md5V.\1
// @>T))@0JGQCH6.Z]DOH,R\H6FW5IWUE-OP-;\H7GME)TCF@/(2W_]>VK4-R-de^=
// &c&CO1_,):GPDNKK/WGeO<E4DOB=a,MTZ#:MY2DTWE]4)T6-Z?,Z.(e](1<dIFeD
// N^>WNf]Y89F(NXX<9Va\^ScXFJda<-W_.)77EcWT@X?9.2A1bDO1V14N/XP/=\Nb
// /<Wb;eL^IFMU7;c8.KM532/(:G2eB/#FZ_cF.?/#b]eA=UF95H)585HMY_3,,CeY
// C+#MZPY:+E^R6O+Qc=5V6FSB6WYF-E74_Ed,eA89gW]9d[d]9N99^S6IL^G[UO9)
// U@>8-9#Pe/Vd21GURQ:CJ+3_81):H+GXIS6:S^#E</T\MbL41PVRHg=54CN;3?>B
// KYNER?D?#_=LX-.\);0Y6YQG(1/MeQ1TZF)]ZN44CI[FI],7G@cLU7).,gPUP5QL
// F<BbE+05YCR.7?&58dYaQ/cT<V+J?-^?+A3A>F[IfAP2fe22-SSXJ=8BV2@9[QZf
// R[H?;SfFHZ1(>1(0[I\FQX490K>7Y4SaWg;1?Yf=NF\SI.VdCgEVZ871Le;#2<@4
// LJC&-^G)S7eQdW3GDJ-La&\Z)5&/G&e#<0f6bbM:D6(a=?E=Q>F8A=@EP32B1AL/
// 7f&TMZZ-Q)()YV75V)]8A(@939gI&6^T5CfLbe+J&e09^E0b^=X)a8f&cMR1>B7[
// +#2.D]?V(;/W?ET\Q;Y))KXM.M2=MW.[7H09BA^QFE^Nf?H2ed^+DS9f6;YTM#5^
// YL8g&F:+K7,@8AJW>MAdN4GKZbff<1,+(ACAFBJHYBV?Dd?5cf)-W[/geaM)7Qb-
// GT._&@>9KOHJYeK(C3KIO/;Q\^HeeF_G?5+Ic8Q)f?M=/_=/?&4<&6]3UN+#0gc?
// 5I\UY,>6\##M]YRg:TPF,X)6<0IE\UdcZQ9?Qc=PWJS>S\2ff:R08YHKVSOaUPfP
// #_A\<Be_P2LB@U0Hg33;PFR&(-)J;]S>9cIQ9T3:MUGd3SO>cQ;LK0aLIJ(L)a,]
// Z^.>S#McL9.H3]07Gc=)6:GO2QIG<7DOKdgIOTa-eFE0AeLcS5HJ9K/2@^D]UQ(J
// DM^(RAM3CBBEM9caZ&IW)b/\QA7#4:8ZB1)2gN3BYSE^g_YYR0]U+0\6+2UXQ6IR
// INL7c6gL1CMTa0/fY;4U4&2M-/\deHY^G5,YV4\#g7SBK[.VSFbM.R?DC;B>bDE@
// LS-?SQA,N6<gTKLA@SH3LZd/fEB]fT(8&8FA1=D^VATIAL3Y^5)<a7#(JK]NK.L^
// 1X=WHL.C8:BfX#dgBNFA7FJcUGGZ(L\Ug+67;]CE?U1STBMRONDf/K=TEJ,U:a_#
// IP]aI>F+E:>2N(U@e1,ZNPGLJc.G--g-F^>V;U9c8bbOM3V:<RY<gU8fM#N@a::/
// 8IBSHe#1f?]=5(4_J:/92#&6fgb#9^SQG/E8^X2]CU=BA2@gaXXgRS?Pe@?=cO9[
// bLJQcQe6+@LWFZAKEcN,#2Z]/8:9F)d7-??SI(\g6c\3bXWEO2O<IG-Z<WOJC6Nb
// )-NUfb2cMK)__LP5;^3G^2LU-:_d\-_N,ARdVgB#P?cKV-Q1F\Z(Kb?E\5OU&6JV
// OL.4@MFSEMV3&X=-X);OYDX:#=TG2Kc27[OUd_272>\\\:3.gJNL?_41Vc-0gNN+
// _3UCUCRDL<S?R;Mb/bR._5^Ef6EN5)C0?Y9JML^S]AQ:B+1gJYS4,(I\G&,;O_BA
// 9].)Yf1;gXb4P&1_23@Xf@9AI2CbW\_,[&9Ufcg5@Ng=)GD60EYDTWS]40B&[g,=
// ?X<2L6&CfH_a.P=b2@B.;J^OdCL_D>@PJ-@)KDfAQG>-FKDcY6=g(aI=;WZ1_d/D
// Jc&MM#^/5&8657QcG30G\V0EN9JKJTV=:R2+>GNO?EZAY?UXCgSJbFJ[Y+&3-PP7
// 5c)dUM[G48]V93VK\T4FP+.He)3P#f]C#]9@d)>VG/]]RUd[dV<=\d5V7A,Red;]
// \aeLeDX)P#5UC72D(g&9)J\,#T=b73U&c,-TMW,Y\;H(:T/YIF-166eQ(Ie2bUCg
// 1#)C0D(<Q]+L:#0PQ:BKNc2-R[X,6bBK/fUA.3Z=EKB/8=7\#f_--166WY2TWC57
// KX3TE2__)VG/WGA&5),#Y0=,,0RMQ-J?e0@5Q;:F24#G0cZV(?d/gN3d+Y2W(EJB
// 80^AYbFLR/4FH598B;/]d<R2_eC)b3[GLGfTS;YARgG[T4X/VTgIWc3#9,C-WMV&
// g(O..XP6\J>ZH]L3@DfX8436@a(VQgeT_[F:8__&(XJ_H59F&aC#+9?FLW7:M0A3
// I-4FO;g&3GM;+a4N]I(Z4W(gdQ8JfGXC:.P&0ITUKgO55d^EJS5P1\0&IT8P5^dG
// LBQC.SXM0Z9S1>]AMg6EfR>FG=+.88=d(dKRAXDCXa7aE?.H4<T77Ve&eEbOQBJN
// Y78BA>WaVX2DTc2464aCeIC:F[D]K:=E7B#4>Z]CREDNcE\L.@K;@GG2UKYL=e5=
// NCUDa]&(fDW51Y13ML2O9K9d5Y)RHFX)?15N&/N[0A3=>.D[94]I,EG(ET-a?FZ:
// A0PYD4g7D[)Pb?BRg\H,bXS9f@;V:/@6fNW129_C_?TUId9.-8;HUf)ZPWe,XK+f
// B2e6JSeI@[NT[aJ9A+]\9)\5LdJg/RIK<MV].L7-GTaBO[&.Y-H_Z&]Z9+XO6G@+
// )BKaBV9=c((V8^/_>>>7E:>D^[\/I66PCfR=6>bA,8H[6]WD4MTDgJ;-#Z.R,c@L
// Y(HFF(KF2d3F9bWQ:.8Y3F_A^7CTdePWD0Lf/#>ecW-;a[<=Z0:EEIeeUbV(I2\S
// TY;d=X-0+B@FO)(O_=\:N&729LT#=)7P)])102-eO];eI@ULb0H3<ZC<[R4bf_1S
// :5#dc3<K-^;2+3[O8QKTb-LR<OM(=IJ.gQG1V)eeS^B5C/)_3,+TZb^dQ-12?X3O
// )Dba1G&b3(2YDOEe/HfJGQUMf7;]<b(;4M/>-A&M;W;^96G^N#:-?Q7Q:)MDHcg,
// 8[^d:K^TUd7&Tg(?dGS6^]O/Bf:8V[Y/^ZHQ6U).JBbEdC2#/]VIH^2S--(Va+;<
// Eb^I(YHPSffL85GR#MF,cPOSKT[OHNB)g#0;F03.B4dHd:R^4[dX4I;1cW0A9\ZQ
// =7e;gGT9ZZ,L#d4:c.g))>:S_E^GK:MfN0?-KG<T.=/-A/4<)KWBDFWPb_@\B5WB
// 8Q<=2-PST;2>1ZdFDf>@F<7g_UL@>^.g5NQe0c(1#AaaM>MJE1QM(XSF^HC(PY2X
// Zf]KR8N?/5QN[^A\STI<)DHg]5R7(RA,RXI4L@&^<;@e2#DS2I[7QP2?=L@Z]a#f
// L?>gL)FTdgE3;HEKO>WbJ_eBPc,\e#93]44-d;<Q35=59F:b1=a.gX)W:5QEdOeW
// R7E[F2Z7g?WIg<cM01XV]L&R7T]:&AbCf]d+TCEHU\1b\+6&Q)(e;[6bRKI-BIW7
// J/Q>?.22GX-T3_OGO4G34aU4>KU=X,QW5c,K).Y-PPXb#cX9H8(PKWTQ?Y>^]^gc
// #,\3,,R0+7L(R2F(_95UCb=3?W+^_VIKJZeAG8MGY-e;NWJ\1UC-^,D?P,L9Q89C
// -,XO&^XC)<03ZHX[>_TL5G]QRWI\(g4/KTDf?;?Pf:U.9dD@R,=6-60W=OJ\\FG7
// 1=:d+5PJ_7S;cZ3(9+XUZ0@DJ_A7#>S1S9)e8PWE/cHQKK6_L(/0g[0_>,7QBA9>
// 2HB605#>eN-)GF+0e,5-RHf1KUC[(\>?P):KVE3_^._^Pb(:6E_SRJGPOYQ5B03g
// I>Q9R&@Q><bcD#BF:IcLX@-Y0B?.bDd9UDf./Gg?5IJ@QJHg#WSMVRP^.d]a5VeU
// /\1\WaB5MP/eS3[B[2gNS81d;M;e9W]EF=fO,f@M7G>9V^,3]^-gaP0.S&EH_X9#
// 2ff.TD)[+8UA#I,W5\[?VWbeT3679=\&T+W6<1(^FF,K69Qe9_0WV0+<U5+Oa7PH
// SPT4Q7AbV2(3GN1_46(,/WFP7K_d)+<KQg8c6->OQgJG,1&,V8Q4]^IK#IG)RcOd
// \DH69UZ\J(,Y<VH1Y]gG2,MU#6O#+A9L6)YOb;K_Jf^BaTI(235K2G.YO^1c#3?G
// G#ZcI-KRM4LP/Pa-HC7I#X&QBaEb3@_L+++e]G-2L\G([RC>Y=@+36H233O(5/2W
// DJ.D>3791Cbd+>0DRWb]VI(eL+Q+Z0SMa(?NLQ9XIEDB^V/[P#0I\^#-cOb;#\5d
// ([2g^C5[Se^F@QQ)YB?b\(CDWTCN2S7&&Q8@PBESSB4/7,K0fNe-,/99GZL+W<&6
// a=4]K\gC4)&ZaI#R^Vb245);-dPJ3MP?+R0TI)-Oe.fNb&SD3T)U(P.B_F>_(\@&
// ]F/OSN8(&UZDOWe7+4#VM/CI\0dgME9Of5ARc\<Tf2gL+?/3;1+V?(IS+0N]99^(
// g?4Z@[\<;]Qdd4/UEM4@M\1)^?@<&<(&>9]REGE&#@EccCX=9-ZE2]X4P;NYPT@5
// ^TS?6gd1U\]=)H_dAXPLBM7X)CJGB2A.5@YF-7cP^ZF<(CPTeL:AX8;C[?TPJ:)(
// 2&T5eQb1YQUUP^4+AR#a8)HN0UVNG8ac,=[GU=aB(DP9V+ca;PPR4,-&WaJXDBCY
// ;FgN&KC4Ze^9L,_dea9Qbg@)Z0XHOd#_]@)?7OO1?SV#PG>8B?c,MaL:JGfSQ3-;
// J7E<[((G8_89O.=2B0aXJJ8BHC\3_CT]QJF)E[/C_O=A(CT8CBXZ&M&fY33>^aXK
// @X3+FVNG1_J8MP_:Q[?)DC/SYH9#]SRGW]5e-I>>e-\19M[TP9/@\GDbb^V]8Y?#
// Nf_LdXeOSRfK,[X5[0DV1+_=c3U]Z^D)599XAHC?V]Ea:;\H^<2C:2gJ#-R]b=DO
// 5EPYKYO<L.9;.5[MB29aZS>7a<.ZcW\[=^UQc5b]Lc_dMP192DH8cd4O:/(QO6&9
// dLK#>,]T]acJ/(YZ;F;,BI;#FIAAK1&6[ZJEfZB3TZQC:KX?EZQS+a<79S,6+&EW
// 72IDLE4@e@Df:T+2I.d-/SYG:^536UBB@G6B6+CBHW4K[#Q,Q[<^2__I(<DE]IH(
// fJCJ.3HcXf:X/?/KGGc9F5FALJ[@,?VI7+<P&YEFLU,.Mc5CPZVRacHJc.T1_B(1
// <>2]I#Na9X4ROcYT]:8]1MfeU^#RTA[HNDVLQT+,?D;ZT@L]c,2e/CDLe(N41=cK
// cVb,BJVQ>[R8SOC)g1GBaaY<_Y3\,@.9fBYH6^4EJEH/EX;^6,5J3RJ&gCA-V7L5
// 7&RV5Y>gX85R>\)S>S&9.G</#Od[[@?C6cJQ][E2N,MOgd7PJLS\[=G4BBQGX\L5
// X(:1BGBR;AHaT(Y6V([R-9V:PB)5Y&@-cSNCCWY=cWM343b^[gQ]V[b.I&1UK.Tg
// 4NM>(L^D=&dH@-_aT,^cG@CJM]5M]A^4U?P:[CB^6@F_QaSIVdQXZfIG=;=\X@dD
// 1T_dBI-678U6Z/1PV.DBJb\aN@6>J@L1HU[6-)MPR,3IW_ZM1;?bZY)./a&5(:UZ
// <C6E\_:2BMPDV//GCMeE,,T:[]#/C?Rf<<3]eT01BE<f-/e8IRZY>SP,a#=(ZQAJ
// :(X&;TG1(_bUXL+))d=VJZA7;dX)/ML^8U)<NM81JNI)a_OO(?(fNV&U+P35D4))
// (LPS]R6AMd]eXd\a@AB&=(@Fb<WHVAEf,9)#\(Yg8FF/^aM4B54;#2PKG,?eG_6O
// Yb.0N:QTOYT4e\#T/6382b+HB[PXL4/NW@H@;J-DdBX0JVeNeSdHHVOMF=N<LD3I
// d.B1+_10d?H.TCR.WB-Pg53\Kb7QP4)7R@M._DAJ=Z0gO7R[^3:e3fAN3@;eA-E?
// J)>HKC1GgBU=SXH1a<^gXLab@@2HcXMV:M=@T1dT>g,)?BW?8:.9Rc7-G@:1+J6(
// +7d-W&-K])-dGHVY0DM&Ob+NGcV=CY4F4.<JN<-db->^M/.E(9DBW8=P5gSIUSRR
// UJ9XO\(\FgVVP#]V@Ug\G;<@FbH&bS/cUO4[-2G(6(A/0S]S<TH]1QTdaR<U1DVG
// ;2@:D#bcT<97e83].YQDb[RRYKBX,XRDGGYQ4&MC(b,S3QT+d_ea@@(Y=0HaPW5F
// 7G3=>>M:&]05WSRG+D3YZ4DYG+Ke)bDQ>F5,/O5-/K+5>Y([GH7)MG69e0Qb]5NW
// [LR/Ng9;HA7=7<_I<.Wg]<PQfZK#Xc+&7R=7M2\baC54,5eRREWg/TPFe:P.8N/]
// ST_CF2K;fDQ#Q#FLJ>5^<9G8B6>:[[W0X8=]S7cCIfdd]T-P9R&(X7BU1SPT=94-
// Ba3V/KSc6KE/+\>]9^?UG4(UEPOeM=[b1bSUQW3,@afJLIR-g:&1#=P7f3;Q7Hg9
// ;6DXfXAKT9gfLKHTga._bERR.<#@G5:@[U<gER8-D(L<b;ca\ZO\UYeU-</ZeS6#
// WaGbd:82(+VZ/ZI7VB=]NVAQ;-Vf.19O;Ic6K^7EBY,U74+38-.g<#37RV5.IF2_
// 3&#2-S)4HE9M<>]QYB-WH_[.+<T3=#EEaMTY9/;?HD)PKWGN>VM_aRFJVc;&-=OM
// UUcTfUSXTC+S/PcaXE6fFNeO+g?(3Q:&,V+V5_F[/SBUYTY8&.RXY-X:DI:B7gWa
// MMb,N;/AgdN;Nb[@TUOBf[4d@I:09HX8==<M)R;5WD<IM\P&EFe57#[?K@Ie_TE(
// VX\e?FLS,TB;L<J230B7=.J7R9Ob2Y.50^#GF@M.e6A,3O;G)=1+@UR=4NT,:@^F
// YaQ;]_#T3E1K9?I>dZU#?gYX31O\A./>UQ/eY<Cgaba/GO2P](eM-)Y@CT,_:C:f
// N31d_-ZD@/1,NNY32FCM.G0]W^,_+6<I7H,HUb\1aY2DE&(A0f+2)6>=7M5OZ2Dg
// \&FZ,1d@GXZZV[c;cFeb0WH[MFgX;5Ra(9Ibc7HV_V9GYK6T-]f3[_e6H;<7QA:W
// PS:c.)#CP<;A36gJZ.-)Lgg3A48BWJCcRJdH#L\f&2cSc0>f=PIa05R@U,;^McY5
// LIW[f@&-.QUTS@A-+EF5>D8DVO\SY3bI+49=\JA-+D#ZT9=1E(NL\[U^^XX15)I7
// ee#aWE4J32bFD=ZUf&XS:LOE)]9Kfa;(3a7B[LTE;ESDKGf,FX^65K+PA@cD&GY]
// &N7UF-#gW=(B5d3)Jf7/@Wg>S&aQAU>J[gM=H(PB^4TW_b24_4)Y-CBYB>:V#Q6Q
// P_KIMR4U?cC&LXH.LK(8\T;Re;,TZE,2UH>2c20&?1J;4:S)0J2+eHC<U7Xe&1AK
// P[-Z0eg2&-9O5YK)EBd,.\)+K(R(#aH6V3AKH,L/+/@W-a<?CD_)D#@_JAaX9HX#
// b]PX?(O2ecdf6E-7;;g&>CLQYVSK(d9&S3_K]Kfc4E4#?0eX\\>NTSW0e_=^@T&/
// QX-)YE&a&1L&1\1caZ@C0O(,HbLf7X_6Y[WL0,Ac>S?]VDQBPP\NODFN)7M@gd-I
// NHM/Qb&&0[a1PgF+2+V@X?)f1:?1ZK>#,B:9-178gW6SNH[Q\_622:b8?6D4WAcf
// T>CY3DETb>8SN:?[JK4&fdC>:9=Y/c1#d6H?CFC]OLcX3_@6A;HY:6Yg=W>38c66
// 1Y1,E_P12J\3+L3Q5BJaLe/\Nd8eHT)W\7^.N4/Y@_9G<&&2fbYbgS3bQ]=7)D=+
// OFL+K#PeQAdUT@fRB4+gK7B\)Q[,\SOCQ[@\L+.3d/:J93eWXK:4+g4FI^56?M/g
// ,5U:f?42O,X?EX;KP_,E8/VQTC)\_;R=eZ@-\?A&cbH(NfI4Bg[VZC7H0CSf++O)
// )DK72=5LG=#EA/4RfYGVZ&=OHIX13?VNQddAAJBUA1>C?QAQO:69[_eE4D]WMTD6
// A,47,07Bb(cD=1-03Ke?,a5f7<b1D;5c6DN];V4.R3SHAUZ^&6O-cXB;<X#()]e+
// T^9DL:GgH>^>cZ-Rg59;1:(IX(TDT:21_8)^[^H6<L,d8dVAQ547<\GIBGS(>F5a
// 7(YRNbKB7[>e-^1OF1bRaJI-ADCBYE3e)g2QRP,\,04#N8_BacPZWT?WZP&fc<a5
// KOG9]b]/d<K#\AZ/Gb<Fc-82:C]XaY8K&cJ@NC+[K00>,KK1MNA5/1]c/)e)8=@d
// EG2Ye[8aKdB26g\F&(EZ)0O<IT;=f-Hc6N:)8]3QE+ebXCAf152gXDTRPcW2PC+e
// -[A7P7ZA-V=G4Y(EQISC_I#0;=WK-#CJ(Q7eI&C4KL)QV^W\KG7?@N87SJK=^5(:
// 8E\.K#?g#2O5\+P00ZGXHI_g[E<02XL[^A@4-[G11/MFd>6J>G[GOC.4QGUYB7Ra
// U38c->W,#?7<.C5G1[I(+FeV_YbdNHa.@;U^]YH8=adOF,+SXBIQIO,>8@&1UVLB
// d7ZE(2cA:XCcSgU77<.:V;afJ^Y:Ia=8aUaZM[_Y@:FK4,+<N/:^_:85DVadZTU9
// F0(+23fPC<1gI=UPMB6g2S[JcXVV^73R\VA6/D([?SXV]#e,9_<>1V.)PNLD8J5^
// 29BMV@D?08?ZY4-_b#/fGgHQ5bLVC0#Yg_(C#N<BEI=?(J#eJZbfZV.ZOQZ./FT(
// K](K1^@&_X8Z)TMCEG<_CRfeg&_gYgYP0>.);dSd5]H_[DFA^M7AgegSCd:e:d[N
// NZBBTaLSMCFU1_&L80b0FdNM_A^CP/1CYW.-]>deO_ecBE#K[O<FVI+/VUG]b&3@
// ?VO]---<C-LJ?VWdbBKV2O]gBH,N(Gf0,.[#QQg[#8N9W(Gd40dbM?LQ1M4/a@;9
// 81MIXY+UO&gB(0D^Y,FUJ3AX3?3RAC18?B9e5Deb0/g@_>)P+QR3+(KBEN7Ve#@&
// AKK60>\H=M[>U:7._\75ZcE3B(Vfc3N7@BI7=<@<2PI2(P_e9C/AFL4NXa9Z(+1<
// 56VOS8fZAJCL2A<D.X,VfLOIB1IR&:OQ7V+[AdAKXVT^C#_?fb-E;DaX9#:H?A,V
// T90[DVKH:>@CALO5^VR&GXN6UR]\?d13)+(E?dT]PAC;F<Z4c,>47ZM?.C5_=C3F
// e98YT^R5D6Jg:f<V58+#)fA]ZMaZA/><>UZbGKUD5Q4M,IgdGXDK[&Q5]J@FV40S
// dE:,b,=@e.TJa(6,_Gec>8=#/PZ\\&#3.Yb:+JE;5_Y(23RT+A/MC)(#?)O-ED4L
// WCAQN)8A9TaVC-&LH5K3.37S#dV>cFaP1Z65N=994<b-ReHL_/P[?,Ab[D50f9_<
// SQI-D+V<a\PFaYJ7?IgGZ@M1WPQO/0(&/W(L<&TJ;+BWR8UBd+-f7J3?:8Nf<3Ad
// <S_^[I](Y9A97WY94Yb67bdH3J/147/&Lg<ZZC/B3Z7:@:Sa_1b/17]FS.gZ^?Ra
// EW=[abOCEN)P<M3WP_/<c=CW@EXbL7#;ca1=\eaQ\5FALNZa64ET7+&M@K]ZI,f4
// (>8_=KdC][W0\=T.@=OeX5e.+(8USSI+1U^3<bKP[XQ)W<5^(HVXf#8H)BU=,T?+
// cdZ2=cWF9H6b77=L;G7H44Pe;]H7VC)T3)9U>:f+CPVXMXOd=VG8-+cf(AP];7IP
// 3ZK#>>,O-9J_<N:4R@+W0\P]S:DY)eWRd<7EV4BE?,IZagMUa]a0\6E/H4J(d,VO
// Z>fRK6R\H7;D4RNO:Z>QBNV]#WC>J[7H=cWIfSW)J7a,/@fTe6bFYa9\.5AWCP+F
// g8#1;<)(39@6]J9V87K0CVQD4VGHeP-Z#b.+)9g]B?[EN#bYXZ[XceQ1gVD9-HaR
// ?g0=?dUS,1DIXA#)+UI@<LD>Z7c-Y0:W#KL^_+HJgB_4Z.5#[20BX[UM8-/UU7a>
// /bD4&T6IN?B</IS3SUb&.->2\H.46><KN=V)AV6>^,<.2Z:\:Y:)(182a,@[M79N
// AL]<[[2/I,,]2?..&GE?N-cdW4Ec^?9EKRBJ,O[8Q+FfT@SMI\1eS^A=16aGaIYO
// ]>ZPD0#5HFX8-&d?62A3Jd7[5N2V:>3I/9BBST.577HE3T4#J&c&Cf,57L]S5+^Z
// /G-BM+L(3H-?Te.5]]1Z&dR\SDE)?W3N;.VZf^576S_2M]BFP5->c(FH33=&1S@3
// 7,0eC5FEL[&CE[EI(C6XIeAeXP]<5a-JCZUCS>3S1]LbJQ=SQ^I(LTSC824Eg)_U
// +Y?XHDUGM4E18BdQU_dV^-=T<9bBgRZg_X]2FMc2)Dd85L0[b&UG\CSc>8N2;ET]
// g\M0&/#7:CW)WX^.X)-#9-B;ZZ-c;MSTCHb+QeR\_VZ&YPgb[A>6-JKN[7V9X.3[
// F@&51#9_OP)Z4)>C2:SdAKQGG\^A+Q0M,:BT_I,M:XbC.Q@WIeO+gZQ+b<g^#EQ:
// ^GKDI>=Kea;UXPEcT.Te;6d=2E825e;+T,]#fCN?EDX4_Z5+^QML)5Kc#0,P)F,@
// @)F9b=gWD60L^004W,GR6e7Aa7(cW.W./YI#NNY[@f).><:De+-?NY?J@@/gXSMB
// fP40MIR.4/Q.QZg_:50=E8DDcVB8GTFOa(M+La)MA_c+R2NALII8-5=NWBHJMM[9
// .73+eK\?V]eQY@J>M[&Y#M&\U.&Y>Gf7b+8;Ec-5KRg^PP.g73J_].?2Me;CCL,S
// VPe,0BM,8(]QDTVG41F>a#9.4)P?g)H&-UXX<fNJD3O.69Pc)[cALY6]J9?>e6[:
// ,LO8W)Y&8.+.HS1Wd_E_dQ^C[XRW4DP5BMN&2e1<d+>:Bdc@(04C.,bH(g]K63@f
// 7]VfDcKR\Y^,GOfYGI/Q]1EZ@Lf7SJO,IZ:&6XURFe?-_=W\PXbAJU4[=&dAZD?4
// R3A>c>Yf,eR?=V)bbHgCcY&-g688G,>,(-WPb5\+PQ)+LD5LZ.\PdSE_2H.BGCK^
// 8F\:O[;Te+D#/f:SL9O)e)O9IPHL\.eWY4=?;GJ#?[8[dJ]IZ(S+)VTG4LTNbcF+
// L0_dH6#eJ3(Q=:HaMSXK-b=N@X(<Y,9UW>/JRUaF[(;(OAd[Xe,6,XYZ1I,>/(]B
// aY2)f9+VWUV?/>BI6>BP:NH]BZ6]I/DV7:KX[7&5FV0;g,4BHOgeWX_eUE5RUc^(
// 61=U0:;.YK?/DXS(L4Z2H4C02&Z]c3Ze@[;GR2Q\0?Rd==?OZ)XWZGT/4+DH=AE(
// &e6;CZV/7C<?QP,gK)g^]ANLQF(2\@V\,6I9g]2&>gY_ZSRa6KD+N]16R1]X3fVA
// X1J(M&57gP@1[(9=40XV@CHA]>VU6IW;ObWG=H_Q6&.CYUJ-dONB)IWHFRb.=.a6
// [;.5;L4HfY/ObZ=/H?;^@8CRB1E]PF?JH1[=6VZK_YH:?[&VHAWW0:[UeIPba3;Y
// cKS\&dTRfAFA@(2.b=4,K=Cb^@(SgFVVMMCQ+YPdQICcg)/>R<R1N&JK9d3c]Z:B
// M>7@,QT/KdGK0O&R5Df?B_GFg.AYaVL>+0V.M^bNY\)2Cdc6QTBgF-B_VNQ+d\(&
// WGCg/HX9MWA9QDE79a7HWeRG6+GN\b8K3#VN^-C.4&NEf2^+&M30,D)RIg)C_(Jg
// _5g43W#FQ\\[5(L0R5QI(83A9KO&2C[e4Ib]g9-KC0fR&G/eS)_aPJ5)K/S<0:#(
// /RE;[g?=eA+/Bc,]&F-VXL8[/U-;,S\3aIY\-;6IcI9_c:f5B7>Fe/05121)95EP
// .5e:5[SZ\?)CJ,?P4?]+;3&YP;aQ[@AC-3[CF_2YVM,KL=:WI@g33@@gTVEb3+@E
// [)eF@#BHGYe7>gP7L;DLgF9aJF0-.9[7;]8b^+[_7I>aTDX)\Y(KUF+77cHY-M\,
// a]+;9IEZVO<5#AfSWO\a/ONUXQMd4FYgW/?;/.&RX.-::Z.7_LWaVQ7L@e(^N&6g
// =gD6[Kf16d9JCJ)3)g.@IA0,Q[ca]QC6b]\F&C/a5]1;Qf7XB7ZS4&-ERdAYK)RQ
// N)3-QO&JZ0#HMWHC2?T<FW)BE;7e8#MIR115>NM+bdec?]cGI/?8a/eB\ZWD<R.b
// VH?MP(T&:<Lc@8f3<QO>/:#]?PSY,U1_M<g>Y0-128>:eK-7c=W>>\<e08@CA/MZ
// ;8)UZ_+U)CJf67W0=)40?T;899,N?UFgd2@,-0DGBA-LN2f)SgAXC(bULL]/:]Z0
// 0/Og&-dZdU6X3Y76L\@Wf,9FX3SCWSY=M^XE2+4FT8S&;7@\EJ3QRRV];Ug);)Bf
// 3/:Q>0R>J4^)#5/0325\ZN:FZ3&7b++P81J8RcC:1.4@03][Cd<II&S6006)b\&b
// ?O<9(CU8F[FKaQ,07cgf0_=TH9IBOC?7H,&TYO77N.8D@BHF_Za-/GcJE9FKV6Zc
// (gcW42SZU=KP560P6DT-VJeV/CX>#>^TGD+>aLP.Z;g+]<A4LeNg)9G7B>Z:;VQJ
// 9cPE(8KR8eU#/HgHN](YI/XV<W[XQYA@+:+:(CeJJL1/X\TOUIFLN<N)[.Jd9V1.
// e??-)e-N)NM7E)-4SC\XD@b4<1B]S01A?^ESba0EHc=([MSBb;OAe@##4^;#)ZS0
// TaW&5QGMe1?;JI99cIBDVA-OC.,3g)^:?)#2LP0(.gcN(+gV?L()[G2W@.S&/1b=
// 21X2CNFG&;ggEd3X0I(O6VNOC-AbZ;ZLZYS.PA],R./^=KMG&#0W0J-E7\R5>NQb
// X9.]5eZc-6F([^+_&=L(L,&bJ><&IJ2N1EO&<K0/YLRL/)D^TE+b^P\[Wg:M:cMX
// Q)QQ@GF48B^_^PcXfA4,WNB#<bAS4e:AbYBe5eVKMU[F]aW?5><\HE.5W8;W49^N
// QE(O\8E0;4/+H@D[bRHR;)>.-YNLSONCZ&LN_SaG;T?)U^/_>=ZM0@M8Ja]DDPW9
// JBA>^,370gP&6JMObW?EINZB#Mb.81QYfa5,QD>\fOI8Fd_=ea;a@b3V,5a-LG=F
// <[0R3]R1&IN(F69@eR\cK9(SC^6bP+F[2)HD,EQF7#^4\\XR?+5K8H=?Y=T[H>_M
// N;ga?8GX0-==?9F@e&H?2HWT.YIB8<Z&a8LZ1_^_UNT>5Y,4:/WE55>HFcV@])MV
// .7P88BK4]-#AW\;ag+CK<AV9X#fGBO=O]N(-WJX];>9JN/8V7eS3S8;TR)R=e5A(
// >:K<CZc)fcZOf-^NO&g8U:gdb]VdUB(1gR9B;#3.c>GZ0ACfc38RbEK>d#fXC1ge
// (,+aCL<M>LD2bUC@77@0CMRUa<.(-=5:MYJ-@)e+8F@P_K[63EY&DFF6/&dcN7Wf
// \+f?9K>2MZ[_:UM>c&7KI3bA29geg8J@FGV+?S3gUYT+.bR9+?LGCP.)S,HfJb:&
// H-Q4Jg@<]\^\gN37RV8[47GR<-W\A+^PPO,f8W@B<5dN2_e8K#Q2U#b+?g22H5XK
// ae(Y,UANe=ea/;bBM1aR7I9Y^H3,.NbYA2^KRdHK4S732/>&S>;FC8)0Z6F_-/S+
// 19FZ35@aYId15g@;[a+#^ZGBV(OD#TRY<7LSeR)>@<.[+-,PU+ZGM-4^XYOJIK;V
// aQ)3P8CNf@T9=]>FHeOD_2c#M[F;2)VPF2e.E]/_[RMDWXI;:+[KFZ7g\8FXf9H.
// PS7=cY078]O4&QP&K2T?>]PEKFQE^PI@d5TUZE],1(g98A@0CC\M0LH5=D:Y&VX0
// <IW?_K-Ed;XbF;CBP<OGA+T<1MOE(d3_^T?3KLaWa/7]^5a8>dU4Y5Z.LM25B9;+
// 3cf>/g+I#6QD4c/J4?/K;K]aXKI&O^^</d0V/FQW>J8+-/>EG]F5V3+=^Z.]GHOK
// OeD+6J@&1S4Xc,933L=LSLS>W(bR2KPW3_1S#MSP4F\TO7[+\bXST8/,5&bX0BG4
// ?HeQ\,I7+AJI+Pb[;^\GT.8V5cHY(7,^,b]\K&4DaAK:A>fcJ)CZZf>&B;/DJ7_f
// /,NbC@+I+d<a07MSgC^GW^,0@5CZ4W<ITI&O[QFOaAN6aYA+e&UEPN([EZ(/AGg]
// >KH;_RP)^24DZY2SaZ,XS9NX8\GYJ&5LKI\@:(RJ-)L8D+S8(I30X?.A?)XX=,SU
// &7@4)B#<O39V:=0>RJSUK\G_J/f__KMIQP?5Sf#+<CB5Wg9R)O<E=267RSJRACJg
// (e9YQBR)O23&FT#dK7fG]Y8S/XQ@b0e@UU(cSEU/:3VGS;RgG7?f)_bJ?ANRD_MJ
// ]<W,];XA.=:D,V;3>dc1^SLb5ABW3NVH->XM#45=9-G3,fW48QCaRTIHXMSEQTOC
// a7D9@cJ3b<F=PEfdYWb7,B,<5+/F>V2>M[]:RAJ;H)M6G#I9)acbd)USC>DXH<Y+
// TN6J625Pce?7>X5@KKR6(SASLZ1dJUSMO;^@C\aA6X/-18HJ@5SW09J0:JHTV#\M
// OQ3)IKFf1Z,a,8WN4L\^QG@Z^;C2E.c@UA<[.eGJe0^F9S9TE#BRK(W)-#]g7DK>
// g)B^GTDI==_A4U=5#[+4_e=.6>0B0TN(FfVL,BS9:5LbTU?=G2/fB:#&_H5REX[:
// -TV?+f5K,gV]4PRa\^e(X5J-QJ;VVXXAGH;GY?2_YU:-/8F6,EC-Y]X<gQ<KW;Ag
// .cMBWZ=+IV5.DI/g9T:L^Ha#Tf5<6/G?[P+Z9d7e:RGG0P;1@WcG5&8>3+b[NTX)
// ./OLcfWX7/GI_&A7\(7X\+U:325W-Y&cBM#Ad/^K463g(a[d-b0V;TJC(Jgc_E4C
// D[Y?gYN+c<Y;8M.8O[DcJ(GTOKN5RQF6b1:/O<Xbd\6L4+(<LFN@cB(=1KXB/?[1
// @.+@L?NCX8MTd2XD^8=2<+OSIdMe3(#eCE:b(LGBM>[A4_>#+BVgEG-@g.5\<Z-<
// d6cBS\W>/eg,8Z)eH;Z2(5B(&UBY#?).XP1@7[TSMaf<PIKcPJ00KQY\gSa+M4dN
// U1IO&^A./B0U<1AA,Z>@.0WSfW:4QO(&96c.)&I6#;\K8VKL@-;R@>ZY+03+1BTC
// bHR[5@J(fS[:?0W+PR+N(e6(CC[HGSD/#RaQ\#PfaC]+;;MU;P_#ZE4ZWNYZ7>UY
// Q45_bcfYQgS&O>HW[Q<P^d[^c<Yc;6,W)dOI17BaDPg-8Z+B-5a_Gd.TS29aG0P2
// ecYU2M[YJ&aZP^8cO2OW#0#d_X@>[O/bN[<^UN9G-<5)5c^CC_@Q>8cC+YL>5S>#
// >(<^L::04GfCS(K()GfEZ>&R]9T&W@S&6UXe6BF_-6TK&Og<</5TV4QMAWc-6H.H
// 9VY=51+;N;9&_)b0#a(#d=Ka/;27.8Yf)1[d;.&]:;VPFSN5>=-#ERb7J_.,2?1?
// K:aG3R=&MXeZKD>Uf:PgAE;3?_2=GW_gO.+#f<[D,U/B+E94_3@JIZ;<GYdbd)S+
// C(Q.Ve?RG,.e^IZ8:13TSZ(d-.dSN::45\\]f#:8?X4AfMH5_?L#/7(>5],5?4]G
// Q3fXW8JF\/3Z&L[^7IEaTSK<?)f@;;a/C&Q_BE\P&@,9#:L]G(F;@XQ[^O=57M0b
// V1?#7Tg0=H]WN@N903HPa_cTB4P([QKQD]J+Kb)\Xba(>#f>b@Z_Yd9)>FZ3D3J>
// 5eCgEVJXcf:R#]DP+^WM^Z\+4cS@CEYG]=\CGT2@(Gc,N?]6cWW)2[6CfeC3dQTJ
// PFR:gKL8GRQ]3c;)\>_9)^d]bCWZN#UEY,O<O4;_#FB2A[C1NAZB1A&KNVOfD236
// cZ@PF#,D(^ag3C8YV7BY3KB\6F=95A4NcW5eQ)T\54M:GJ7g?&fZ>ZV->De:L[2N
// R(g,V0T35aR@-WLf9JVR]\5gCg8^-1;:7TJ+_^5a,&Ja.#)\\CCZEa0S2._LS,<.
// ffAE,7WGbVb:>f0Z0XEU/f]7bcCI8QFY&B.Y^KB;V?dWFc.b31+EI7[M^;G_Kc0D
// <5YPYGM[3-C5<A)G17bgUK0Jf)ZLRST9;S1TaSZfT@)a)1TcF@^_CC[1e6@T7?a1
// 0IBf(fU/U09UKH,9FNeTdVA7,+HX:4TbAX,9FY.@3)V;J.(,\N9RF-RE(H75<=MO
// 1GZXf.ZVXXHdR.J&6]K3TF<)6?I7SOB(+A/O2T^fb>-Da,(@IFa5K#6A>:W1S,-(
// JWVN6>OPB7UN;-0H/.aRB9_4g5CU?f>#]bHVOHdXXBVY9;0VGS_(P5VV0X5Z11Ye
// 0-fE]9]a#6a.89(QT8K,FC-[c][4/&9+>EBC]BeSR)-(MSB+7&?A;)M@U7D3OTEX
// _<)9MF^aCdb5>cR#IGUCS9Rg80/((:=E3L/U]cKF;M,d2W6Gbd0a=V8ETCRA6LWg
// D?bc[C_FT)0[=#<RBe?dQaL<.fA?_BYNc+:aWVU/CM+^Xb3C.-B#OVF-]9GDZPS_
// )gBaFVGGMXNAA-Fa\.YGC+7(C7MG5.^cWYLRRNY&27ee5EXW:YEcfZ<+EJSM+W7g
// 052+,MHX(HDJ^LZe+>_D1b-3A[4#VI^c5@7?@@_AI3IHTd0bH2>.1B&258NLXe,K
// OgFeO>8-L_#CI2adDPKaE5BN,:ZG[ScUU\=+e@F6[)LI&SIbUV:f?9\eZDEb3UMU
// H/&;aC._1bSWS;3;_[+9H&34(K8]1N]]&GNH6/B:>/WBG[c8>M)a54U;_)/5V:Eb
// ,KL>4dcG>>8gNXcg?f&DY2HPBE]@C?TUde[6T^A:VD1FR=LgQ5@_da@eHI)1d_SK
// D^LR2KgP5YAE=K-NJ,J]2_-#V^5)d+NID=/:aS@@?JNOA[1WdAO=VVc4DSIL[Xgb
// bNb;#.0<I7^b<?+FP=RA@7VQaPBR2C#6+#PWK)T2R/]:=L.+1eb#4.A_L+faeHC6
// OAIaJHe1gH.1F/=W;f#WU\B?c(9-/JI#5O=Ae@BaNId8/,ZGM4(XdFAc:dPYCOE]
// R_-4TcO)8>Wd#VVcTB=D[]@-&6P;+4D#4-C^U5#QQDg]Gd6/L\J))41(M4Z5Yd:U
// #9467QcE@O[D;[FI0W34)X]fDT(T:0SUKOOe9:T&+KIb5W+:^^_5QEEg58>_Y.^U
// O[cCW(cD7d1K^>51gE(VOcg[)&HcZMJ7>&;XaQbA9S9a/0S]AU/a5K4RLI@D)-EQ
// &0QSTULI@CLUK&)[6+GV7dTY2WcB-dIVA_#BVR0[-T/T2a;g0HT\Z27S.,1=014J
// 6ZGN^#DMN]0DCB;beccNd([P(^^gPGd/N,?5WA0>(H&e[=O_T7N[Y;F\5_8QcDV#
// H_ZZ0:bAWY:0OR=0RdRLOSN8@LP[g/P+4NH=+UCKe]-FcQOM/:5f@8TURA;UC6P,
// GFCdEb<I>0.8?f&Q@8]<8A45cKMf^ePLX[U_08P]UgEEPOTZO&-[TE&F49d21d13
// 6M]FJGIaAH:]g>-2P1WfX<]JQ&<N.dQ/YZLT\2F[:\C<,JYR7]X_V=W:b&c1VK0F
// F8_47(<JaVKEC(Cb&5525#(68G),E)-EA@U[H5S-A^<S&]Q>d1c3R^D4]@X8VZV2
// Mg5#aO5K;U>afV1YX/96M,\)O[S8@S5??6SO\cC[0-fegULCVT;Neg\<+DN,S<gW
// S6E<&,Yf2EIL#DFW\JT)-D]21Z\214-\S#ecIE9&CTe,M<D&6#._bN94:c)gg1O]
// X)JKZ&3)A/Ba@:?+d2XCe^\O5VVbSFO2^bMVGbAcf&M/?1/8[C\Y3S;?<^V<(U3,
// <_DTB._G8];\_]YTG(W)gASN4Sd3eJV+R4.;)R[\U;)5I5IfQ&=(=UNM9Rc^=;#;
// ._Q<Z<(aU5N,NO59S+AJ^6J_<8bX<J;^cJQOQ)@>=K,-cS?W+O4SICEU@DZ[0<bg
// U3U=C3O?NE788&:XR0TE[WFM3.NR?Rc@-g):QgXOc7B#K4@K+6+>FUCGSMX^aT,;
// EQ_X(RTB.GY6IB].5T:>7>+-O5JUDG=-Y0D#b5Dc3G5^_+->YfN<;UHJ75WR65IP
// B;c:&#MaK\:X9RYa6dHQ#7&=JJF_6]0Laf=&N@VD:6:aKD0>&VgM<Jb[]T5NNCQ4
// DVO<]XSTE99a6(8?GI8(9f?Ea/#Q?J7D;&<)3QK/@B1IJa#gcf;PMTYRgJEf0VL(
// U;(g(K4M,QA?.?9a\-O#]T3(31Vb+0f;dP=C)XQDg-4U_([Ke:611fb]^?T^S<H,
// aNcVa#Y3E+ge;[^IWXT[CM?W;(X#?WC[FU@)J6//1XgY[K^L0NG+2#DW5>5f14:K
// +_()=dEf.9a#RE\-&=fU\)TK=A:&.E8TdG+5HW8aQ6VE)&^&](\ZP+,)[KI/ZG,8
// g>)J:UDF:HdE3(SG+8_)0&[49&3BHNg#]]\K\5M[_5ZRc;U9a<Q/[]H/SCgVMS4V
// 5gI3.5@?=PI(X35f6dIX&ZYA]1da53F8\#ODVOKcO>@0FcLcZL.0-7DI:UX.J76C
// HB<D[^0_7X,U>c\0.2eG<2SUb>/,&LOf7:ef@4FUQ)\fP[IS3&=Z=Y/2.V64M@#>
// KVRY[3c)f933A-W;g2J4(8FB:?,.,C;NGOaCJLWAc^cQQNWBR4]NX.)gV=&(b@=B
// :)\d@+HNVMHSE:[#bc:LC3@fVff)..3&<D?WM\^N7JgFZBV#fGb7)7\=VW_)_O4A
// :aEK]([RF&]e.ST)PAg6g(U?3=d=g1NAFeK#)88G[@<@F0HeW(YIR/N6965.Q)gX
// ._57_dA,D;3&0I,6=PT]W_2H_8[;J&GaA+:9ESU,W7_c&.QP9eD</E#T=MR(-)/@
// aDb:Y]9Q@O#c2VMBMRP&?JS2DZ0J^Z?^ZBf4NV0d]NO?[&>#X^-4#(O(beWFAMKI
// C5D7R()ANf<Q1I]7/4Q3c[/5V?.LfYc,W01A.ND#0JDIW0FZPF-G66#DEZM]7P+;
// S+UBgfE60TSea#U69;YR9O&HL6UFH^eKe?IHVa7^aI+c21Z[ca198L)VW=8(J[G(
// 4];HX-a\&W,-dRS>gK##TSDNX9e2#Y\/U.F1W[,WL=OWN[2=V:gPJ10cC),IK&UL
// SbfQ,S];F#_3;K<e;,9=NVA:E,@(;)_NE23D#GJ[PB6_8?f1BY3/JUeVWR)V,GG(
// DAK:872\T8G9&Z^XTJ@NDP7J3Y9U@03H3dWgV=.OIP.eHTK_Y<g-V8dWNEc)6W-.
// N7cG19bZC-J_c<CK40V1YdLfMb+5B;E,6YARH2FBd3BdgLN;P=NEcOWWGTA)RYK5
// Sgf=(WA-BBFN&=T\<f[0P?5/W#U.W77eJH[.d6fD-V(+.^SPV8CeOW&1S?AS[65^
// KObd2:G@)FD)=0@H:-F??9PT/T#?<)_O5e[.35EDTY3RC>^UI[;;_AcH2f-HO/UJ
// [9e^3@a,P/\5f(cW&6[1Qf.8<cXQ6^<42RMRPHWC:-N(2JJX+c66ab?H6^18_?79
// BC#KaXJLV#.^ZTDI2SIPR?/5VIF35[1/H-968B/BP2=J48SJ_2A;(LLT0CC_WT0P
// NQ43?5^a0YaQ#)9&_XU#=_:4M6;\4@-T;D5BU-+,3Q5M==Ig\KD3_?(E6;Y>.X-)
// TS[[+^JS;\>MZgb=MQaZL3M^HJH2R1V22QN83ReLF99JN^76)7>fSSEb2N78dDeX
// )eG&g\WH#Adf7X+ZK,C#ENe8TZgP6472-]J5f30R6Q2]]4H4V38)_G:ELU0QcgNf
// \=@Q62TBT[/)-D2F?b1.7^XJd>W@.]\(<QSa/d[5Z@2g+HD7BKFDU/^WGQ:KSH,U
// P_R#de&e=V7S\aV&AN;IH0ZgUBJE?ALgV6eRb_B]BDWWWWKXPK3WO1Y=XQ+=dAOI
// ZfL,208.J[\YLO2eb)-Eg1;+2U&U?SJWE8IcaI4#Q?0UEaG=?gGA4D:M69cS?OS:
// FgLIZF(#Dd7Zc\MV_,_bf[BR)A1XF;=3^X\8Gf6FK?N_;?_#__H?;Rf;PJYID73a
// @P+R-(d@=B&P7BTA&JPaO2P7_NVafd(-PLU,9N7]VM#/UD/52J:PNP5S9aZQYJSO
// M2(G,[-WgDea^S)T9+e/9U=)UGXfU;PSWZ]00d?YPH8+S,daY5a=6+NJWQeC)=_P
// c.ZZHa+CB0BQRY8F73+90G@V/K[&NA:_agb&.EeXZQRJ:Sa1.8AVZ=O,@dd\\XTc
// D@3Q92A#c8V7a?0P8]dB-NA2Z4GebI:c;b<CD(c?Dc4N<2V>F68TZFS(-96F6Vb&
// D&8Kd@WN]aV/C#eQ#Uf,S8]KZ3dJ+Ye..UKK/gQZ109WQ+>R[T_K.cS<AJII40cW
// Z?,@bR9>,0gQ69TQV5f@0/V^M1LdeKS;2e&1bRgEA\MMYZ>,4GK?,J>TE^4SK2U4
// BaF8g9],Yf\7GHHdWA<0?X8Y8Q(3aZN762#(NEGCL#PWJJL25#Bb;V^\E>LF?PKd
// dDcQ.fNa7^81,T#[b3N]e<:V^##bbBaT4=BQ2^()L_R@f9P&g,ZB>e(4dX=6/_M6
// 86O0IVSJVMSUOKGTFS1TYa\HMX:3?X6H=7E/UW<I>ePVF8D1+5fR?4Ced]b@UJ(;
// a?XYE,?O=QZI-Kd0JT.0?F5MNE&bO40]6Y?4Xb+L-7[JZ;DZL(fE7\MEPO?GK2)Q
// :^1BFI/W2R^K^S&CT.dRLW<Td6W38?O1F(VD;B?_TIIfX6H=I7f8BW-4d7&D8?<P
// @]YKT@^6P<A[ASdM-#Q//&W:&S1B4]71/_IIM.UM05e929L2IJ9@W+R[B>B+M-?U
// DXe[aP/dSXF>E).X/_Mc9DKH:]S.3a.M257.8L)?PfgbDTA/NZD&ZEM-)DQgU.@2
// ]cM/U_d<6,<8)YB[[>BQX7Sb>;/7=B[2K^X3KfX,Gd6+.U<;&&F0(,#,1>,OL2\D
// S2N6\U2R=>;Q+U5NKaUg;)2JVc-1@8T\MY=gcIfD+g[Pa:b.DZ^;.(@+3H;:RI,8
// <SCBbD?3X6_IFgP/eY#?<2N4\CU/d6W)d,<3Lg_OE7V<,cUdM)d:\X+=cRTCT?6+
// 2H=8(+6FFTE7c/:c#d+cHfRO\VU1VV(?YY5G#WHE3@2[gTeG(g1<Y\cL;7_M8VIW
// <[O6HW5YATUf^3(eeRDDg1MM^8b>:FcZJM^C;\QPGHPMK,\TN0Wg;.d1L83^X4Ud
// Y7JS/SY+<&:#eb9Xc.U7g[,G41;<ZL#WUDb^]/PY^17/@:E5cH5@@aUe@VPc&)M1
// cXMW<)]?bbE)&34-WJ&3c^VZd559YVOJ>SM7TQgE+(0,K[JJ]:_T=EM-5:L&0\&g
// CV1fUX2dfFZWM4HB/B;SgfJ^J7-:#7N1eX^#55_D.N]H^K2OL7;-75Y^=aP<_7d^
// (4E>+I&dQP#P_K1=J8UX5Y&P8JddLf]8XHc-M9-NMKKL6D_<7F4C+4Z_?US,8KEA
// AB;-)>_MKK#]NYe)gYNXc2PTa/c8][1c&+\3,L75:(=<UK;JC3M[G+FIYKL6F(0&
// ,X;]c]M-(1:4D.RXEA?GOKKBG96eL(+-e,O@#,.1=W=4&a1BB_Z36V.4TfX=Ug[]
// P^_45>H4ZCW?,76EMZ7(A1S=;>Ld#BXd2[1W#YBBA[?9[:KeDZ.N]ZSN5?dU1#D+
// N<0\gV_(3=c&-4f&dD0PS>gM&;9HE>X:H\N?^R1(DLI4HX]21K:GJLd[Y>68K0-P
// 4-EfW9^N8B<73O\)\J14Y-KTTL/QAS-IfPBM=5=N=ffCGN(fDLg9HX(/>ZBLd85D
// E=O;N?0#?dTR[eHcX+D-R>9DQRaS61\DJC1,N+,OJ]b\,I[Jg<^F9fH0:8>3gb4+
// O=)2BLXYKC];1=5MF8db[c6XONK^ab-564J2Q+X5g^)-#7[259]9N6KdQgeQFF<2
// >g.,d]6:?]/FGeTDTRVR8[++^bS-U0)A.6&2P[0>Cd:/__\]A8GW;YD)X2fH7C33
// U0X9+Xc6+,?^2/M&CPM6ELKM;D).8IG2AQYB0#+4gB.;1H)Ja@S03c<HB.LBcW_>
// GZ36_Lc-NfS4WOSCNW]Hg@9UD&CJPc?MVaAgX_IKV,1APSYYRN3faE7KdXYHX&NU
// /#,37:Nb2E5b^RcB^,/>L^W.S@)(/<_/5&8&.4F_??WQ#TQ_d0f3S]X+Ta[BFD.f
// 2V&6Q)7U5?d/+g&KaXBUbZ5.+N7>9=8\^3+-1B2e@)02,bLJ^)547G:7E.#?<Uc1
// XRFY&ee:\UX+:5cgI=^\^Z(BS5EOFG&aI#D93DQ.JR:,N\>MC6C:BN][(UX[9W@d
// N<K?LA3aUTCGb4U87+2C,:8.A5C:++IO)7)-SE7;8e=&Ff?b.C6-)3aTK,[a\AD,
// 1.SBC1JV]TGbS.U9f/MAZ\U4UMLB,Cf-a-@YZ@Z5CF_96fO7(K#=L3JM^]4IN^=M
// 3fc[VN,J^b+DJ=g,.7D;1I&YDfO)VJKe_5OPde2@CQ>;#EWD4MW@c.OBgg(H#1M6
// B;W56W_M+bW6]P3KS7I,N7W]5;8a#e871VL#2P77H(TKZVag6F+0J8WH3_6+_g;C
// c]WZ7T+93AD@.QVGY)?^=DSSQF6UXZ7REU#KXT/@#ZA;M>=]7XCbAI^a_]FV=R>5
// PKHN0db:/9Sf[HZOC:a58L](0a^-@?/#3@,9TT#7b0cNcROHN2CVY(B;e7-aB6V^
// f8HM?Y18+4ETP^^-)-@[F88G:3=B)6H?XgbVOPT(-8:R)Ne7)OWU\6#Q<@,ZKWG3
// &-03@Jc/B\R+d<0\O(9PE36HJGC18LMeRL8FfXIA__=0CT0NX:f;LRT3;9-QJON>
// aI3UITTA4PfZ[.eJS]SCT=O\XXH[VTgI(7<7HXAHJF#)Yd[A>]a:4&S<[fWWb>gY
// J7:QVSE1I7G^RO/E(,KLT(-Yc1TL?5d[J]#bES&@0Z)Y8QKT#Y3g=6WbNEY]M[0N
// XG9VU=J^6<>&\F+M4T_2G&Aa2.^R\JJI;g[=CZBZeV2<-&L_A,^fV0fYB,6:fT&2
// J,P)VZe)KEZb<-IT?X)XC]K#I\b32SOWS+O+=@b8eHH48A+1b)8BJZV_F+6bYRVS
// )C/P@K]@V=fdJ)59D;cL,#KZ&dV.WUNU_<:++73_e\0;N4D@A3UbW\RJSgT5[=?2
// ;1&3TC@.01f4W4V&MY]&K=1TOM3a2@0PAS&MQ90J:W(&RZ=(Z2Q\JP7HG/YX7AB2
// G2/0R:^40#0#PZR[a_SF&V:cG8:>1=CK:08D\5J\REf<g<Z5M@H<AHdgSG2M/)9A
// PD[J5@B#)L+ZM.L?-?(be,>T@]_(bc+][\fIV1-R5JD>HJ7bf].9cNcXNJ@L?2>&
// >3SZ1-#/K+7F;Rg0ZWU<Y+,_^]+E/2]>]MV+>&OV-TbR8/(5UWdEI]NH6ed1VAL8
// aIbJ?[CQBTN(;eVC:df^>R6I&2/K]aA=],/MF_=F?[]F__9Eb#3I8[5UP;eF>a+C
// 06FJGCJgSgE0EPFBTGOQ>U[6c;5,65249@;O\[F2K<NcPAe;G7O?.b-eO,2JP[HT
// d@\RB3J_FWFc5S=645WFWgf#MC-U&:<J?/B(UT)LB-=D716_=7UXeK)(8/P0XRaE
// =;3&EU]4O2\@RV.]5>KIC/XW;MP^PH3H,X=K#E)(/+W=WL[1+S9+;+ID0^(3b<8V
// SHc[U/YA[HVDR?Y0U0],+F.@2HB-SdE]EX(,T;A=Q)NC4YCee/W.b-YQ-_eJ<0Vb
// /W#b<b6Ndc#;S=RQ(?3BPe&(D)NQ,#M,]4C+a+aM_21U=G#C9d[Ye+2]Fa>4+V1Y
// ?DKG-K45Q4d?8HdA8^8)_\;TM]DME^T8T\T]g(F>@c_73;.QMP-@-J((N4F#<B-5
// dR)+4G_:c\dN+^A1a1[L,5&M-R,0&S\138b0,3?K=Aa()a/UR&#<#_d?c;VRUIEI
// D?g@0AUJM0&YECCcS&CEMaW8D=,9WXPJ#^/CKG4=Q><ZQLbY;bMKB31fH^T(09#K
// c76dL9WMBL6,F,.61=>8]8SGT3<7bGCQQ?18)bZa7R3ggac;=&MIP>+fa[NBAK:S
// _c/.eVU=,fAKENSUBYc#?7W3Z_MB7HX-2^d4aFfC+I[RBFL=H3;H;9&WJaM#[5->
// 7)9&gf@0P@,/.0IU_NIA9HH<]J.aefDXd5JIf+R+CEG&DO^D@QV_abEG=.f#K^ZN
// R,OaJ0\93;MFSE7909A+KZ<&;+A67eND-,4@d8JV,=EL1f[2:1\D.H1+/a/YO-E(
// 1,3dBAW4cTb.N8CgG@9,&6MK[c#g6b\5]:L#;0,D=@V:OU/@JCe+ZDM4@J8dEcaU
// 3&0G4EBdd3.4FF/9g.-ge)c,bdOH6O+:bfJg\\d@eZ@?.ARSJ@Sf@Pf@fYY]&\^-
// 83WNA2V1Y8ZIg-f6]+\V-L0HP+G#\eQ8fYJZ8bOc82Z/?8PVO^/A.>f)eGBK78@[
// 7^cLa8]R\LSd1caP2_b.A,<]LcZR30PHMYV,aa0g\fPVY@<&\,3#1.[]UO]]D+Fe
// O;6<WPV]@EN(U\6K<X7gF2Pd8]E7,JK1EGBJ.^1=V2TTgRC3a[a^f][8],P@\L^G
// KHc<=C=Ec3#?_B80ZbCE3B7D/F9;-ZP=]1gfM@gDB=de^E&80E#<^H<H.XY],bK_
// 0Sc2)gC\3cZc?9SUSU9?.=Z#+C&JGBUe3I?ag_X\;78defd<QL)]LG9GS@.T.PEe
// 5D_B.KDBDO,8HYT>SL0[LC>T=+D]fdS3=d+2a]2811NEX<Y)EB/([G#R^I(<#3Z]
// 17Ld^/G>23>YK#>(Q=_KN(D<e2WYeg=(=3V:+G@>941MZ=?>3)ONJFga#O(ZM3A2
// 42+gN6QE;,P-Y/YBLb[9=:R,P\=K;ae&OF+I>eT93K?T(#2S<EUU+XaE0@^JF78g
// &Vf:_;A2T4WAagNf=J[E2+d+)9]df]PLNOgI19a-Jc&^XGYKQM9#:)4@dOMAF]WS
// A/7K:RPD:BO3D9T6Y6.1?(d@g3DU8\[g:&#6)eOVXQUU-PZ=4BM..]UC6[Zc4\>f
// aR1:<>/HXTT^ZT.eJ,5W):J>GFSM]Lc.0fCN]D=6d]0cP9^8fffHfYCb@=,#BK#g
// IeR<c3J-BL:K]b_3KT/dPc;XV8A\3[fQ(/SS7E/5b=A^<,9[Y?DB+&>^b:@)2KI/
// #R2;VX;EbH/;4OBIf5dd0V\8>2M#KU441Ge8V\F=Va#8V8C#+A_b\#g&\D,32M:7
// M0YGRfV#a6I5/@@=BM9-KbU9(O=Z/]7/YScM?VCQ\ZeFcMe^-XS]NMCT]8NVHS+F
// OKBWe9^Ee7-^-@d5_HKW+6KG(:A)Y=BIO;Wg55ObK_CKK12P=9MAY<4G(OQU1T&Q
// =>>=K25>KaNI>2[J]ZZgA^;9If^LN472fG7)HOB-PUQLMUaNYKP9d&O#KEV7//5]
// XM[#W7Pe01NZ.9fJbJW5QI-5b1-eeZFMFY5gMKC<H+O+R&KQ3T>d+)gQ1D?B6,a_
// AR,W+&?X&TVd^KH@T+\c);;Dc^/-G:/5HG:)E79;K=EX.3aCV--_Jf9OW;D-XMc)
// Ac0Z9d&9Z9<b<UE9fZ8V,Bf9Q4#]UR3Q7O4V>67E]@c5EH1;7YG#?:\-J#^ETd#a
// P@E+O<I]WYIB.?910FW@X7W2R2:;,LO60GMEUbKLXRcLX\G@7=#SG;6KeCPX7Q@]
// Xa&[Id5F>WVUf9W(<d(.<F8JM?.f?38MFS_?-S63(NLRgSP)3R\R,KgUgTg#:A,&
// AA^R3](8>FL\AUVK,WS#,FJ,A.0<,(PF))?c,)R>EVdeV/,JbK4H8D)I1RaS:Sfd
// ;8,37>JUGIWR_E67#C6&4YSO=dDGNZGaTa/B0P5A>;400M:9PZ;gZ[VG\_>E(6cQ
// H[MU/ZL/+cO_X-8,/cV_d?GXK</\-88Yb\KLCM,_9#Z/8Z)+gEVIg<W+<WOL1<:-
// @WN)WfRcO6g@.17J<+S9MRR8N1TA=)M3W)OHQE[,6O&d]9a(HL;MYG9DMPe7:H/<
// @VZT_9cg8A^77I53@BH+>BZJI4/1.ARL+AaDdBIJd135@6_:5CMZ7A5X/316\=N7
// 1;R^Y_Y3g_V3K7Wbg)4UC3MDg,;-NVNce:,/=@VFFCOGBX/CX^DCFU:0U^O]/fMF
// /Y@>4]OX\(Q?FZMQL06H7;O4X]NFJ.?2+6F8RHg5>=bE9S^FZPdWK,&=12Z8A?K+
// E0WX(U?(dDQ#L[8B/K9X0AKIDQ=OZ(>gbHY18LAM\=JaZe31b1&097\+WEUS;d4M
// \de6^:_dX:6GZ#URE7BN..>8gK1;;81=\&.gec-OaUCWI63;HQ<&1M_[XSI&FdVS
// ];C4?K:@VfDR_A&f/I8Y#+dTX[<EVSX(M=^Z@/Q54B7T=Ab0?.K=G?aaH&eX0b,(
// 8#ACP,O-b5c@D&5]2A)R<c;e,4B+Z+]R+F1aWCT;X7Kg@=]VUNK3@Yg\2Vc23^MZ
// /&O\9B9T/A1\C<D\&#R94(6:E(^H?C8@#ZZ&M&)UbBZ)D99#CKO<>XM&9X48CF64
// :5HgV7A#U@PA/-bc<]Yb4>,V]d+CZ]dY2c?(&.ZYFZW9f8CX3R\[U3_a42G0_HWI
// gH)2ga9c&-H[NY0<()^3ae-A1,Q<JTc/V<g[;SY4-H;A=93+TMU/X#2;A[J&f4K^
// PDbKUXU0AL47,UN+A.HWD>ReYT^::]J\&F6:BU@OPTU;cf4,\O&)>:8IKBYd([(V
// +?>IMSJ0XD-XW[L\QM^VL9GBUW]3Ka:fA:OEF@74fBGJB+g[ZGB(BQMJSL=AgPS#
// SGXcL->ZMXGXLV/a,d^@R+d,F,f8HJ#PJV2gP=AN/f@+_XT\[(HEL^(4)H]M(,3[
// ^H@D@6F[&U<fU>daP4NGDHDRJJ9TQ^b/./TQ#B#N8J:c<AKJ,_2I;XDeVd0Q>HdT
// ,\#0ZYPNFH-gcVCg-PU4,./R\RR2]09gXG?d3M2b9aVFZRZ1UfY>?FgMc0GbC\BX
// Sd.QF:92;=/?U9/IX9Q-9;M_K:ZBc1J5U0FZea]<)fQPFd34MUE9bF.K(]ALI_]2
// ?UZI[BAK5Oe\4^4LANM&e52X)5+(d4bWBBc:977g8cGZJNMJ[S;R;EY\QVDS]W>Y
// (4e:8B78WKa[;6.W6Z[cbHS>?O<861FD>.M>>W3.@\I5+Bg2,):F_2?]aQcYd.F&
// >4He>-3L=G)dQd]P4e[0ZSB_SORPaK2_eg;dZKML;>5Cd\]S0JdXfSKf,7;;@?fe
// 5PVg/#:+K^OILMDdJM/E7QPB?X];dZXWWX0\c2HgfgEB9V:T<TE+;,7JK#<+YFL=
// #C[e=P)PLYLWG:+]\ZJ^?&W2aER9-2S=-_NGA/R^KUL1]O@Od4SZF@0fAMT;a#K0
// V=H9>2(S:ZT-<ScgBL>&f=K>?aYTV@^D[KJ<.ZF]4V[5faC#d/IJEgaV(]8/<-RA
// 0B1Y9JIR>eX_J1-4^&Df>O/CQ1B?E\K8\=+GeCPVZALe7VCGfXO=&&L<Se#+BAWf
// C5&8RC1A?d3?aLZ<K,[HIY#OGb:&/:_)ROJ>\M,9SeAOd:;/6dJGM9E>-#<3R]+\
// b/,:Wf@MHf5eY_W670\)4]9Z,@g)ER5O8D=N_&#_Ufe>QgM<fb2J-ESH4e&I.6de
// <5FQgg\LY=/S/fZef7ZVCc1)e6@8)e.=.&)5X3F0UHSE<F@6XF5JbI8O&/C1Y1-J
// #U[X575a<d2IMH?=>TeSHTTN?eP[O<[4:g&c?F&C+e_#29X:dHHB7Rc>1DI5U<&\
// 9gc(<MCef3[f:2TQb8F#-[L:6_7YE)cEQ^1eOE:HI@BL/Z((gP@gX/:6Re2g\S+]
// R6>&4BfSGQ@b4/H\MAG0F<6b7,ffIZ.(07@0HN@6F>RD92fGW.(gBE5M]Wd&&a^H
// L@BCZeRcP^aSA^R/;I,3b(+D[X+_:9c4P=2S@/@8:dIG>.Q?;=4G;N>>>/CRG]HG
// dP=D/U+@;2Z>UD<Bf2S^e\2AMQ47c;ZA1d&UJ64[13#eU&6&Rff@1gUJM4=3I7N0
// 5)1SI25<>(\-QT.4L/H/B]Pe^J]gXBF/DBBL?[5G.<4.>afYF75.U7?Zg.X8R5a@
// 7ARU&XAUX0Ic[-b#DdVZS0GZQI^&S?e.XL8;/>,N6?&,d@9Ra,#7X2XVE.+5>><&
// B\@@B7gFR5[e@KRW1[e=8H_U-,;:eLg3D[G7N-C(97<\]VZTNd@)BT2:<&U#Kb>)
// <cI4BK&4_,,9;O@?=7eC.RGUV>>8--LO<((15(RW)LCN#@:5@\\47#8<b]Ad8-#L
// I._?G>d,\;PR(2PP\KN;DEXCRcdPE)5-_GGX2-A&B+4;P?2G-2a<=1\KgaJ<b<SW
// (K#TF[,g,BL:_:b::1MFM.,,fg9#PT:+1O(3:FJY-V4+HJO,Ob2JL:dL7-8-cf>f
// ]NX8,OO,E[;>+HR<R.[Q+>,.3fX6#KCKegN\^TL0D)QGaG)D7d0-NKY63]B.UR6#
// 8?DANZYMB4M-]CVB2+\BQ\6J=cDQ<QLPCNV?(K2eVHL/5ZDQbW49)FC4K#ETNXg6
// cd++I9JKTP^HX4B/H:5ZBaL25J^T<F>[WM\^>g?1+E[W>SGgV4CCbUC38L^WU8Y&
// RP_(G4RMSQPBI)dRGITceJYSgbg^YgU+NGP=\b(-\1c5,;?2?H,:\+AG85-fNUMU
// g:IBe:4Q_N.fd\-K]OBaXYV:Zd4U:.:QH4Y9Dca\<^4(ANOW,_5cbfDe9QPRI^8E
// 8Hd+D^A6GG\&R+WfKQJY@?](LQQN_Z1<0&V&Z>9f-RUF<L0Jd=cg2#e4E,6?73ae
// cA)AV#/CRJ42?:NFM>AN[,U+M^@M@gP#Q=RBB5P-+[Sd1M6&;=\@aYI&#3J?FbgO
// :SLE^O7UF(=[,?+YCJ=O7(fCA:CNOJ<T[Y2Q5OR9337@OGRRXc.I8_/c,#62N+E#
// :KMa/d-1->G8W@7Wf->6/78[XMZWZ0AD#AG[7.EQ(=Y1)#_-X1:H0(4deERfG=0g
// -8g;_:[<])O6fJ;DSMG@2Z]8EW)R4#TSK3KeBB]]bHCA8FMbNXNM/T0P,+B,ac<N
// f:;T)35b8CPObdU+]],15&SbDd?9?4W&Z/]/Y_,6Z3P?MZ)OaZ^dZ/EMOY0d[/X[
// g-HT00]2/5L:?EOb#1>-;Za0Ga)f>>;M)gb\.H^g2<0eZB27eI/N4SF1)KDEL2LL
// Z[).S3S;4LJ-YMO\C?<QFP4+,Z;&83:3@>87(4JYZUS^MPK_^>JYUPBV1/b6^#?[
// D-eDU8\XV^BMY[/(Q,Q^O\DX[ZB(TG/=gT(8Pd=gD>ce8\K_?KW-HR@=2GKd#fF^
// -)8D8[DSaRB/J7-Y;20Fa=R>e#BSOfe\S81fe2AaDE--Y<T_G^7a#WAgXbK;+\+g
// Y1)\=E21OQG2;e]ZZ<J+>JaBIH8LCC;(B@PR\WFT<SUITFfNPRZCcLABGZMR\J+_
// .LaVgKgCaYbO]<CXYCJ#W]2:J<NX2HaBW0+B2Og&3O;#[#=N+^=90bb0HK9.\,S_
// Ng1_>)>;UXD:8-4d/^LEOIW/75)Z53X;19UGM(#/89X<8#=3=d-UX4T+Y;&/PYRe
// @C\[&]S8B^+(g0eQ6):[PV6XeGL6BA@.T59P,>JRAM\S=XQaebBLH>H^,(L6+B3Q
// >Y^BG_2WVEabZ8<JV&L\7^_]U;0e5EeaRXg1>9+.DbN:1f-LTdP,:(AKe\P,3.I&
// B9C[<[WOg406\-1645P\f90&&WOH0CC;(353a:4#7ZML:XI6)#<=(-7#F+F,]f_d
// Eb4,^g)&)>IA>2G_^Te5)bX5Y,M4TY9=&]O2fP@Sa;S6IcegV@SgXT43&_G_Ad1H
// -[(A_b,c<b(eR(7Fe#eUQE0BfA5&.&3;KH,gKGYe&YG@826+3:<gC[G]:gRQP3MS
// d&][af_C5?64G7?&J.O28,IN1+:9\YKZYD.AJ9FG@1=@7(O03gZ]KM8#TK@.;<TA
// ^+3+dY]BNDAEG@GN@(M)0NWN.BWfT]Y)VdR7T=IgIKX;?ZG?7_eI815RA?D[MTTJ
// KNC)3^IG_Ga_#2b#>@Y5&&>bW:>K4^C44VHAD<8gYGRP?]1BYW&ALML6/KP.+ZD^
// \4I7UOd[,<8^5_A8-H-Z):7X5RRDYY^>-WfUVUc?M9RRMJYbJZ\@.3-7Y+aJW^XT
// EDZA.^_C=R\d??Q/>QaDVeHbcWH[H+NM1K_\1g_->a[3/))^DQbO.6aMN<aQ0.f6
// 2QEQ,V[-N1a(d(QMS)TUOP=1aSg,;bG\O&\VeN0^U<@73CNa:FUL;EI5PVLBHU^8
// G/=Ne8R8V1]T#>0U&eRZ977g]W7#[H^c,QEY<)X?.@-//D></Nc>deS_N#J4MS\&
// GA0EfQ5?.DZDH_UI7dcKX\2DZPLDc/=g?+b:>JB.4X>L_Q=]B5;KA]G02W;5[8Sd
// Eg:dL+7_R\;6I5g&^\H]MP6_g7S\Adg&Vg(1_=B9CNDGO^OT3e)a>-V-M=))GJIP
// Y)1Z\V/AC_fGS.0<bS(;8,28=:OAW&_Z.b4?B5_-.dHJSbA-E:,F6C;5&W66@;M<
// 3_5^f4bS\(PV\aUc,,?bOB9]4GE>]02+DGf](2[UHVVAWQYABW=PVMM_Og<#NYHT
// >E76&]bNS57)S5Q[;.Ld:]+BSG:=R-\[^[^_c:BPO-<UF31c6fN6V2U#O,A3&X+>
// XcWNS4>J/I,VA34]ga.E/?#?0?C-&:1CJ?,NgK;3;#]aDL4.)QY^??63-MJ>7+.X
// aU1ega[_6_Q0\[N-=.-KJFGf2I[P_()8_LB\8_^K]0DfT?9BN[Ag6)BUB3XT:VOZ
// IJA\\a/c)&Ae+D<c5cJ2NK8;;XJ:OJ^ZG9HLQd+]OF1c?SYe^J9IEM(:C856&-aU
// c?M\UgX\G0->ATdN1=^\[OREY\59=fNfCX1<aa?P7,MQC6Q>=2;VW^)@]11eU#>.
// MKcJ_e4EJ@OV8f+^4GPPAM[&C:aaN.eYJT>PRSQ5ZZHUc,(2.R;#?WSd-/,I#,E#
// =O8c,A@125FF=>-Bfa]MY+e\A(_;T<D2PIcC.2D]>SQC=:[^:9=eV\+[8J]FgGB-
// C-7RWU[Ddf96T1D&c?Pf_TK8d]e4IVTL[:RB>@Q(4:;WGFA_MIRAb@14V\>9dN6(
// C-.-7&.S3?D+ZF+@0<1>(F;X;]&VM.&]5,N#JNeaa?>\VeT]ERX-c#cAAW&6DW@0
// W7)1IZ40<5]df(a:ZCf_Z(O5^)V.__[VIY\AD&FW7FW;>BM3XBR=Qf&KG3_c].:R
// VYV.U1/7E=fG(^[Je;OY<g0P=QO3(#V]Zc;c@1LICdb>PDIfN+ES2X9NIfGfeZWE
// P,=-RQ][C.=gO)/5E-OJC(_OK_Q.VdY58ZC\a4A[YM2)((8<g;C]bK.@C#6L4D_W
// #^&]/IOCIeQST^::8bg\f[Z\+ZOINc^MT_d8I)OD1gX75X,^PE2HB_BeUC5X0\F;
// &aT,OYWE#Z5ac\fe5b,A>>F/f:)&K=SE/ObIZ.C9HYcN55-]XH-SFVD^H\,Dd5:L
// 6fT#:g0+[5g+#7C=BX81cR?HSJJ._LdN80[Z4WFRH1:O:D>d7;Z7^4f(+,4cQ<@_
// AC>UQ3D5aKV2R<I#GccJ8(V7Vb5IHS5/XY?Y>V0IG>V&U(A[]QGECYC5,4?]1^),
// a55T7G+bNHgCK1+]E/?[>AZQbH5f1I,G@[/4aXR<DNICffAFD\CW1;1/Zb_SQ:T\
// ?aT?>\a48O,Y=/FGVPG(TgRBDP+#]1V(JW@K(N7A;(Z#RbXGZ;=K=G-Y_^0&&HXL
// Pc#@MZ0J>.JD)3Y,0fSbZ\B<=D8>VDC<+ZL^GeCbN+6L>=)QeJ?4U<MN;JY(eZP=
// &IDSW6514Z3gAR0Zg<@TUS&95+cUfP[LIIb_]/A7HS@2YK)W,e)W0WY;#gGN^fJ5
// R3.\=I<O.9f+:FVB.A);TEC<,Ff&g@[DQW#-/5&UFXTDcACeXWN^[INA/];5:-+/
// (OdXG/6]()<17<3dQ<6\.?]^JP;MSJ#IF#X3f3=G2DJM^_>a)PJ/58DX=/.#aWA.
// 7AI&TYCX<N;,M]eE/;Y(3LB5]e4E5\H/4^@.K(6FV_H9.G\S6IY86f[^OH.@F=]N
// ]C\=C]8SLV;M\f4_M0L0JSMUZ+HHN1@\TL&CI4Sc-g\gL4=L;&e=J-Mg;]\/2fJZ
// g8(gV6+P/Ke<Y/]LOPX\?XX?BG3(&K\ZN8B95T0UJA3:EdMD,b09PY:&-D&5R>?Y
// N(?L_8P2DafC@R:RNe?7F+2@2aX(6eIVJBB49OaN,;PC+19Dd^[e2,HTPa];:9A&
// T#,d-:5G7bH)GAe=ED9H99NP/5]c--M?@H\6G;_AW9K;\,F:4U;e6&:Bg\g,^eg&
// @QFWG:D.,_UaBWDJ77^[e2B@]H2\;+W=8;>V;N-=/:K[,B\_6;cIOgU7.>+O>QYU
// U-E-DTR(@#LI:.2^RIF<@]HR)AAd5@GDK=&?2d,A3X[9WgD,[0FK_eX-C850_^KF
// :fY>,O\bFN^Ee>IGV:?ZEU&)VDS9#B9ZO;L8f\Q#\Z^BSN;/)F^Y0(C?H19,aN6C
// WW>E@cU8,QEX>_8X>;\.>BD<P+GFF@UK\_^dCaH,:8,fQI5(S=JLC-<49,gH7Wbg
// T+[]MA=(W]_a_R<^>Z:2^_@^gR12Vf5aP>cY</]PH0\cg5Qf?HE=>,Y\_NFKMFA4
// WSO&[IHAI=Q2\9Gd@:K.@V?G5C?aT7.A2D]f2;UZ(TU2F#YS&:.becGBBD0^.H]g
// 023/6>db>LFPSPDUQ:bDD&[2WagI[Ba3_g:^+^g68_GIL8\<@Fa6=U[=dVLNC3M2
// ],J_L20_ZT(f?,eWeMFW.S0AX?Fc31;bKZ[Y8=Y#+14+<MUOJB1T=VSg)g=ZJf^&
// Z:f&KM)TF.3MAVSW/D@X.acPa/R;3#;eCWCY+F\,D[[U0HIYVYR1&>9XE&L.,7&N
// 279N;(E#?^(bCM&#1O8,+&MTVa@;,8M0T(\E@@)(..9,T#a17@[I^X[37GP+?>V1
// >PD4[[Y/6I6M6<CTgJNfg/2#ZR@(Tc\cG_6(e[08ecQFb_aG2bMSRU+Q=8[=:7VA
// \M&WJfU[=&2I]W=6U<E389K69+;UM-9g+T:],_9IZMUUDY8-,NW<45D3A^ITEDO3
// 3H]fBT1(_E\:bXKXN4A[)_e5A1;KY@_1<E7@8aFXWQ<+MM)R8^91O32eacPb1@9T
// a&)X\W])._9eG&g4)d7PIT/#Y;OV@bCgE@C9C1QKCB[9O350\@&^5.6,7Ef(GS62
// -4=aa:B3;_D4E-b,]:eWTRYAbPTZffQ6=S?_0aGZ/LW7fPRVFGBBEDOg7@/Z-&IE
// HF2Ug2Aab<AUafa;X22f.9U&362)PLO5J;5^DaJe8GZA,&f8,9U=?)Jb/P]3\b]5
// PWF1X+::9ONO;g;&A<UbDNMJ1/(JD:4UJVC48a@J=cHD]=(#1.WT.I0AFL[dFKO_
// GS7<fUW/BCB-VMC)PI73EgT,^2?,GPCCJ7,0dIMdC_T8_ND3Wa7/[51gIV500(0c
// 6AD@ffcCbO(27TfOPaN8;+b])U,fX3V5C]IfR^.Q\;<&JaB(d6Z\=G&0bb3JVTXQ
// 43@e5\g<WD6Q-FAe6H@@AYY^EH)EFNYN;Q6)E+6?LNCXZ><Y@J^Z<<8f=_Z7a[Z;
// ^a8Eb\-[-=</dTG9#cgI+-UQ>c5(K.D@6SZO]D//2Z36LQKd7TF3JDBK7R<I+@>6
// AEbVYE9e7@X>Y:=DJG+RfHQ=4>1G9gUGHUK4Vf77Y)X?KXB=S3O6g.)fVfZ,GIdT
// b\TC6/W)MV,f:&@T?SZ<<1?aPR)Z3<K@2O+P8B=;[)c,P9(Tf34g@;\3f:^a3N,=
// +L>7(Jc,?<#5-3?/5^1RCgG7M<U=16OZ.)TC\LEJ^L+c<@5^ES)UYCEXEFQ?81+1
// 27WO))++_R(J=S;>P-VZKCE3[EK8c84@]QY>PD><g#:<F?24fX9-33P0+5L+(W8W
// W./EDf.N4MA>_81_2YN/8+gFV[B6dRW2\G3]cIfKIL3-d7/_HDJ82KBC2.<LO_AR
// >F8LYb3K(?AW;=dL#Heb)IcQ8;]EM6<Y56]ZAM6L[&FIP)a#aUB=G/B0TCBd9A9J
// E)LQVC\^.&Hg7fVP=bGS1e)d7/+4Z.G5NOEb,a-6e/2=H.;0W@Kb)RMV.cIY<g\-
// 47gUDcG#[f#M#5gKRW[/@R/cFF]0=bJ7>UL(BNK&1N66c;GIT_&G,6#;#+#=W0+R
// ABER+\Z@fbgF6NFESg07^G4c)PC/@,[G3gGY&&T>56#1KHO#D@0K&UFdHdX8;)/7
// PSQV.3b+?5EFR:/#(ORHS,S\DEX)9[>JZ13#].&5N6C1B9L[6+R96&?UMdLXP8cW
// :#).T2MK12eG.\5@)c-[HX_,]Y:T96BQ;#61cR:VT6eAB=&U4T49N@+a(.N4,a+G
// Ue7#1Kb4e[(K7R]NI03f;WP]\/8,/+BNL7CMdNLNLC,a/4@R>G-K;/6</T8ACNf<
// #VLd1NHJa6e3JYSW,/Ua\?9=]K[aB1)7OaF#FY6HVfXW.#?0@CSP?0I@cHCMd+Ed
// O.fdSBOeE)Tg<V(/23KR?BdT[?>RbOJ@Cb/W[/;+\=Y1R?/-DM_]Z4a_[b?Z=.\d
// 21RJ[fHS6J4\fK9TN@=TLK8B/F#da<b(.e-?OE)]_RK#JET&-+9>29,8QUYAI/X]
// _.T_,H(_/d:7P8F=_fPDP6,OcD@V0+?0X:1)>FN[FXL(/,a[G;E6Q\+XJWF\#/8W
// :GE_D=E5>HT5TA9:[@b,@MV\P\DX;_#f3Z1>JTW0<bY:RY6#4LB.-NaNa(.U0S2=
// dJPR)_1T?R>fb&HK:BGVV9H)P>>3gZS#1J5IdIY86LaMI>4(gGA-<8dV>6SDbZU/
// e6QOKJDfR(Z_EcF>H4e#G-IXA7QW^N64;_9ETXV)7Y-NR[G_.A)IZCN_Q[4V-3?d
// 41/>b1H5();E<^8#(6R(XaU1c9_RfE8F(E>g;&NdOL4a-K&LP5<?G_[>##DZ2B\?
// G>[G5Ne48d0J9#3_/)7d91D0T5bPLR_YW-eX-Y;3gT#2YS)YR1cgd:TBO;(cR[2.
// &_,A(d=B.P?ZH.L,=@ZbeJ20O&=)YMEXDA(9(JGS5:,gG^A,3d;.e_ZYY3,+]Nc?
// \PP?b5TOJ0VeK<KR5(O@TcH.abf0,]?c1c?D.SGVOR<gW.PdK4:HB)Q/-g:A<E^)
// 2@].R7;b:RC1U\_OA1:cM@-/1gF5+2SDd3_4;?Q(e/\(dfP9TYU+6UH@8@H(&342
// ,-9b-RLIg5G1\WF0&\/H&Y)eHRO\1XMB+CY(SZ7\;RE0@W4.+?eAPOHR=gEK@AI+
// -A0+-8_RD+RJNf+?g2a0LXS@dD;3dYfG3/^8QAcKdeJI\2M41e(?,QCXCO^JY?4B
// G;X\=UH5T?GE9SF/_./]]Z0;NQe4-E+20,WVDM00I/[eM8XdfBN9f\8SK9[>Q-9X
// fGb,d;:fdH+@>+>0EJI-Wfb/@,M0X?#/,[\E:JY<S&LS6S2VVMA:cV\)E&E>O-bJ
// 8;?Ue32dFAdaE<dd]fWXR_LA-PcID9U)A=C#N9g]UVeP0gJJ[Ld/=e0Ug82P9YaD
// b,15Cf@]3TbW&I7W49><EINPY[gBD=C/,V+PHdM;WS1N-NRZ5P-;Z[)>Q3GEZ1TD
// 8:UFTY1A8f/)2eZ7\a-]RSW29C@I@-2MB-=g3+AF,K;Z<-<,2&X3dOG2;X;]AE0)
// CX)0:@ZOENC-H_W7#?J._RHQX-cEWbZ;NYU,L3bg=^_BeN+J8]ZSRT2-2/RV5>N[
// =V,_ERRXXT(WM1=eSU/<E[K[=L#Y?BZL<eO2cR5?WW0>:[NK?aVb19QN]8N7(9Z7
// X6Y&K8-d_V,CL,O.;0ZC-N&JW;BA+;PPBOFdCYK0)f<PXFE=f\LQLVE6O4UL(3D@
// E_D^=+\7;dUVK5)B-L+<bD-/3cZFaI]6;KKM0QcR/fDT@\DBU-IUg<U]5KTI[U#O
// N]=.J?E+ACK+U1;HaDcRFR,61S,OZd?<.+(c?&&d1&9;\GNCX]Tc=AV]ID]g5=4c
// 2Z;Ac?eY_RR0dgQK>1gaY3cb6;-P0.TPa+OELG&BW,Y(0Zc\AgGR1NQ6I,=1K8ZI
// Q,B#04VI_TN:]]4&T09J7Pa<\YD#K22MGefb\G:g_:L,2ZTI@0VXLB^4Z9#MV8R<
// 1?QBa+C6YaW,7/dO/P8M3c);[cGX8X01P:KR5J;T?8UW7L9@\JDDS1^Q<J?Gg>DN
// >PN-fB]WQb05A<\Z(0c#.9E3X4Oe]Pg-LVG5=6R+0RWM<X\gBH.&ZB#c12:\c=UD
// )V,R0CID+4c#HB5G(;NM9W>K.eB90T_#UO5b^@NPG+deCa&.VcA=]QX&WD[&,FSe
// (3DgFAbUg<Z6fJb5ePB#bR2dBH.TRLQ&&HZ0g,FU:P8@J/DZRg0>fA69dWC<P1Vf
// +Z,R:G<U/4aEE<ZTJD=V;_O>Q1(UI:7,@H#1+P->H>I4\M70]6D@0.cN:7-]A(6D
// @XVD6B=JH[C3N1<@X.O-9?C)V8DFHEHY7B,e-,R8\e,B=4UX55&>&E1(L9Z:U,LU
// 2;TEf,^#N)58#4_=U2FM3V+0JZPX7@>QR@5BGUFfQZ\T,6S8W/T5=B0JVLO(dg98
// _UX^8K-g,c\_T,fd7)8P+UMTZ\>fIL)a446fC0D[MT3aZ[Ze)RD>+A92.[IKLLAa
// 2G=PAdcG6^fac:&dP&@;&_F?^38;5.BAA_(?\cTXW3J&f5:)gIP-8HGP5I[cUC-P
// BI;J(DQe_N5E_Ad-;BH(._.VP[]c(TJP]1gN>2+N7]6N_MPba5^SJV#aaEB^X=dW
// -PH\6KN\PKAM\<^?1F_NV:OaSSC/B3>BCb(LZBb807c\FF)T;>M9RPSdG+A4@@>d
// ;Z)S::+]S1_Mbe5db>?GTL+7e0cXHTOSTJ,SEP3_(CTJ(RgLS6O,Z3Y4/?1B3fL\
// AdN[+O10GLDR?OW<>dY6OU9SM,\VEdcP,-JeQ/b7f=7?P+T^A6ZNg_^cXdS5HJa.
// gcb+7^A&.=(]\YWQ/e]&GK3dU\N(K.@g@:0Q8&JT)P^d-PFF6e)LR-4F>TaFT@:A
// (&IS,#:3X,JX=b^+0-AbgIB2^HbESI[ZXZ2(I>f@dHXH,LNFAB@-eQ:/a3d5J_[1
// 2GEFFPf]ZOE/F;0RcHQ97+eQFQHJCWDgYCSIYM<AHZZFE<g,Z.0RHL5SRR+.L2EY
// ]8X)>Y6gAZD:KDK-ZMd\^.a,:&J&J^+&#57b5f;\P(C2\#[FOZ85D_U=_HfO:gSe
// PA=[;c<cGgCNfU530=T1:922._8M37Z#)04V\e[W_5BE9<T31XGL/>?GP,E?G;fZ
// PJ^8B&8Hd:aI,XL4?KfFCK#/#0fd))ePT4LKceeIDN]X&.fSX(/5JUAX-7SYD#Rb
// gSJeNI;]dB?F/Lb0/T0_[\WU(PTM5Bf\b8<&H<H.\Z=VRY)<e3ZLZ@(aU3YM)HTY
// ;?+^P5AR-J;9K1<CeWX;;d:+d?eRccRC3a6AP<6eSa8g@(SESY1T\dF(CQ?T?I.)
// (+YE_4EOf,G:I9:H4YV-56=Q)bP:BIW&5d,H.YKC9:?^(191VH4_JNg[\eUE054L
// &(e#-a&Ka=_>aM8@CSER7T=7:ADYKC?O/5XYN(&2E,OOC,4g)P=Z_4OE2S6CHS\;
// a^5-9#2JCK0c&3a/6UEcQ73<HH<IS8\6AZ4BXMOP2^O#/WgEO0KdaU#4d/3+7P8C
// SZ?g91GR6FIU#Y(>be20>8Q,BH:]McIM.Mb^N,cA,7,1P^;]]LaM=2&Q9ddbLgeg
// gIaPe@>;M>-98;aV/IIGb>Q6GK;+PU<I^C>#/:@K_OBA#NYHL)T,ZDE?X?X?F/_C
// :+gI>a?Q=3YJDgH)+D\W53QL[(6P1E-60<^fJ459f2FGB77>+a=Y(42<b+01cY>8
// F8#?TeE7.6]4QQK+K6+d(be8X0ZfLIM^NC.N+/=c:FDKMF30]>AO)^3>:+I3IP+1
// 8EC@#Kf[&X_-]T+TGH?JeY.aZS8D;cZM<SG/f)@5GA\TMJTVX+5FDT,#Z=B<8,.8
// eG&/9H]0/EB1/A=8.SX.YHL#G=7#9<WQUPJD6<EQ;V@abW<[Q>c#2A1US1D([[G2
// IUdBd\).]2^3=&DbfQ/N6gYI=UZfJceYE=&[NcTSa3-HZD-5@.+R;[M6C8;O^Cf0
// (/VP;I4.-;Cg\\dCY-++@P6XOTO/ce1WZCZC9+GPdeVKZB,<eU5\\:FcXgbYTGPe
// TLMC9]<@]KP5+cA@Cd,TE^?ER/JJUJ-UCLG=C3=/J1JY5K6/ZXbc2cFBO==+bg_NT$
// `endprotected




//TA

// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
M-CX5[;(TP#W^@U/J#R4LC@/W0O7GgZ<57D,DG3XD=J>.PT-f^6d-)_49(X]=335
5F,beD2PP@MIUed=1fXTZOZ&a&[G#8fO+N<W+^U5a<9V5,)1@H;]OIeH?eEZaB\b
/d=UD#a_;@?U\H@G9Y_/(>X\?bD1;/g&^5]bII&]NFHdZL;_J>[5eR.29]#:2IZ_
U?DROU;A2<=2+H(Y:gQO0M4G\.[Z4=J>DK8X9g[J-]C1^eH+Z4Z&Q5>&A42O4:cL
/#880;G=+4B/)L/3AcA18-L>P\3cZ&&D+\J#W9<YDdH&^EI&b)M/+?Ge2#@8>S]Q
-aAH3](Q-JUD8b<dTe7P1JS/e?1KeBbK++aGCYS#,>c\#2EG)?fWeCVN15H<A@I:
43,_RePD-A,Te]2?A0Za\U?&W@a<8KaK+4.PB5WVZPEYEOV4(>()/;b.KK1Lf>S3
GIF6ACYF,#gAYC2H\K=VKA&f>)Y,MIK^3KT90gV++De7(cdd&]R?@<b&S)a(c(9L
S<X:SZ3F+Va<G7&;)ZT=3&)gET1,fGS84>OQ2fA+e8aGYI0NZATU/AE<+?N)e10&
L#Z0g7[4>>K/AbC99dXJHU#)PMPH^3Ta?LD>ZPeIFWLQ^)0A481)P+fHDOQ@&g+/
,),+LQ;L0D<]#>SDHP5NXKHIL?+1B71eBeH3RXAN.WC9EITCV\8V[DB/UI@XQBX)
?]Y[#8@7Pe6/3.e+EfPMR-Z8dY5<W<OP\9AQ7?;XgfK\>bb+P2VTGEAM6WNB:E4S
><-/U7K>2LZJZ1Jb8b=Z,1A:J&.b/TAJ:1(I;c;?,<^_<EcQ0#MQH5#f/#AY7gaO
]dc-J:6J]a1:6IfE^K=M>bJ(08XbIJa,-4gSPANEB.E_;d#YU[=O[(6Z9^TM>QYX
Td,7E6QVY66HbK//:=-4BD7MEN=fYF[&5F/G.RY7E(@=eXP0[6L1;4.93E:?Mf6b
,D<gDI::CeP,0b&L4b^?e=IA<_260XGRK26;??#D)A1M;?Mgf?\>+A2K.7KZUXT=
L=WN6X\,<(bTEJ9.[].Hd(G_\FPeFS+QZ-9RXeg2YL+C<W0:-2#5H31HfR?[?+]N
)0PY)PfFJ8g_=FJE<N2Q7KN:aELQ5:_BVSeB39X_4D-C_>1d9,?HUF_W)8[)S16I
Y50]7Yf,]=(324]<<S=#Sf6bDbR]U^g]#9ZP=C^3H:W7gUNfW<bOTBX19-97ac\(
SG[T-gB:TZ20)TdPO8@+bfgZ;>b9Wf]agL;I4:#<T<KY[5R9]DM#Z>;5T[c@:(aS
JX(YRXA:2+)TR24DW3N#7IfY>#H1D]L\XMEVEUF8)eX4]WSI2N<HW^=OB^,6,BH4
_ZQCUcb]D?0NJ)C8a.#)HTKG8LGX3NMa#1_g+WIdJ74Q(3Fg&5?6L4Ig\fR.[AS2
#RT;W[29X+ad<;e8TCIN[.9g<CZUJ&?_BRX[99P=\??c@DCf4J9U1T&VCCL?Pf2M
><>Ab6fJ,b]WbO8Q:g\3d?8=EZLbFdRNf<6<,e,K[CR4G6RPBf/36XPZM_QYGbU1
C3(/D[[GE8f@YMNafYKS1_/T19HR)1-):W6Tb;M^dG_a:AeId0Z(KK9]UL#BR)^M
^H&R9dCRLF-L2/\,La]bE&\MQ8+]X89T^H]]:U_d:W&BQCW<>6)cM]T-\Q+3<]\X
S?/OUPA<.96_]N0&:Bc_Y)\(N[1EOQaQ3<,XEP3XaTf<26J=<N]A>SMN4<N([44Q
/RI&/02=R]J8UV1]9gA19K;9LXV,F)RVEX\,_J?]P@\78>M[MFNDGX69dJ2#B+/(
.?:9:c<>Y=&<;:I]GR_GWWZY.],I08bI2FBDX<6LC_)WP?TYA/M[>FS2U=F9MS]a
11fb)#)^+eW-CHH[Y070>=Q,b<D]UYZ8YJ+b0+g^1acLO(>H]9G];(M0_R9f)gQ]
L)1ea8afEH=<L5\7BZXf?[>Ybed,X>\XabC[8UR&71UE33;#/>5I)/+4C3[bBC@\
Q>M,_gBRTPXTWOVRcXU6XV4NHJ.OQN7c[KNb9:?^c33E(PJBTAIN(DI7D=./3d3X
A\6C/;\cMDP:>ZKI--4DSF(/3-:(J1GUMP:VJ^.Tc8T0L+>cX^PLV?@0O0BL=YUJ
+g2I#[f2V^+F4UYa1@7QXM,NcQ.XEF1gOdEOMFO)Efc19-gdFG_@0D:]EdN(DC5#
L]\?K]EQJA^\\5_5#fe)D2-c^ESOPGY(W_\KJQI5MH8P_DMc>f//6e_c@;V-E<df
ea7-;A_dGM0a\:)CI+IbgHJH6RM:f?g[;1,:aOS.SZT18I3fLg&DO61@;(G6>J\L
W4UG@\(>I.Be-2DV(?ge^D@^M_&JE)g^-7Qd^(;_5UKIJ//LK38+D3RO\\.IATHW
L7=[/8LgRIR1^R71:>>;)@7;\=?+()O1GPFMK)1N-8U5,;@^Cb^0C#3AYL]9YS=:
Z>4U7JF^D8G^3O#;9Ua^,5?Z]PK_gT\34bBN\I63/;D.XEdR9Q2D1RJI;La\,T?)
)9KM0>A8QI)UHC,R3YK8G#GK^<SgL.&IVTcIQM:R&af>1FKO+HG=a=:8:4:b[^H3
G5=2;RN2HB-/C)/de-LJY?f,&,_5b6_8[SAZ\8P;L9f3?_=B:?&[/Z2F7Td.ZU/D
GXb1DdEdXRDD/X)C;/IIR/_]Fe=FBX6C,^P0N8fSHd(/XFA(0&_X]\A;PT./2/-5
<:F_IbFUQ<_R=S+\Z@TU>:dZ,R5P4#)/AgTEI/dbB6[:bKC#:-O4>C^#e/#F,:F,
P/O/adIH<2T]OZe(EFWNY24@KQLeJP=<XEQA?5=>4F#+5SNEgZWDTQS12JIY>]\N
^K<eO@@QN@dPU]K(AET2?NUKH7g1@-:.Z-d,J#YP3>HN4:F#[+6DH(H=>?,Z0Kde
<#5KHgPP?>X3YWM-L_PcKGZ?)1Z3I1[P1c#K:NfIW+EP</UBZEEQ0^e],3HOS4XX
R6cST8E/[_.\1>g&>7U3SL>1XET)c8Y.^1N]W+>TJS=-^AQG3N(A#4)RP#>(Zd-c
.d1F[^4.7SNae=)C42WD0AP1HLEf]EVXO/8,H=T[V?-Q1GYQJ#>e61QKSB=]ZYCT
M#>FU:Ag#W1=3L@eV:Z8ZJ71dTNfA3N5cM9ffc7JB&-2VLMZZQ]=(JY30<5;>c6V
Z5S/<D0M;e:g3>L;g[cH46IDZ5W?G]85HZR_BIccRf);gC_JO5+MW=,=c.+OYKaG
UeH5Rge7(-c]RBNZR(R,2Q(_9(_Q3N3,[cS;4HB&E5L/QA06\[9.9TEMb1Y=S[5B
;-X546K;a[1,?(:AA3?PTB]@D9LH9&6SQ#ca<:2,M+YI0TdOMObU[+]ZZ+>56.d(
;Q\M<VKS/gI,DQ6.I.aTaJ(#4?e2W=KT<ATLgLXR<2O=?V5WI4F+3)-V0;_]U&H+
=CZ;33Y?S:J:P4KUf.fc233GE<ZQK^\a\)<8\I(S]^=9eWe<Y>eVXE3)TcGS:?D_
&)EaJ;eMJZ7WE7YcHW)0,\RAXfW:ScF3E#-K],+B5.:=@>EcH1E]<&<d1BcJDV5W
[Ye&CL28&M.@QWCN<^PTEeV9F1)fIC,Ng/c]&Y5FGG.D^S+.7BI(0AY;+42(]Q7T
-[(RUg&-WS5R0YV(8A1b_S.WP\Y-bDLA]JTe0=E=(RE@X9-U-;-?g.BK@geJ5)(/
ZWIX5U+-PQd/B1=(XU?FTPP:5bHI2ZP1cR+d5R?<VV1cS\JS?=/4&H=?W:e@DfFG
VfLD8@E0&^G2:U&aD7UXeM;)LW&KL&09&1IBMHQ+:)[/W?EVX_+TF;Z&8ZB&0\1W
@e,5c6JOX@9XAW()43aIEJANWGF+FPPe7e?\7W6U1^.SVdGH07Qd#cI:(?2S<H@D
cW1X9L^K?DS9#:V28d,J.M]^]M;GH\7<TSPcDRHO58fQ+6\4;/e22+NBce0F=B;H
<HG&NAH+#P-5e@^eS]Y8;5ZC91[41_a/-=EIWeV;R=VIaSG0<g.601RRK_HWU,e#
Sc5L56KF66P]7a^449RS3.WPMXLD>=-9OP=,01//3&1[-A>KX03NQfYO:aFO^ON-
=GA2GSQZ?^U7W&Vb#0<&F(:-LMPW?CDRN_6D59Ag>EU.M9e4<)@Y(+]L71QLa&#E
D.dcGf(F=2OAGVDc+B[I/K1/4+3Lg4K<:0ICX.\HT22YD<aa13HI@+]HZS._)3ZO
ac#11Q+/#5:9Qd@0+d]32#c0BWR(.HDA6\\?AW)<(Q&69R@?#K7ILL;aT1Sc6>c>
P=O&EN,+ad<TeS86#F;B(R+/#@cg/?X@4cbRcG#a@AW<U_07cVAS2;VbII]-f5I=
A,NMMW:OP/0<\gg0A29=AfO7:M?R5]5=BCa&GH3BN/I0>N7dYfWW>C[^X-;C?5=P
[4e7(.=VVN5U0\BST4=]E+R>#8a,-GZAbAO,TAY^(ESf^:9PQMI84Va3TN68b.:c
[-TE0V66#.=?4,[E6F/(]Hb7=:Hb6_<PF2E\)dF4[?U,MLVL,DYEJ[dEEK0_dRfS
7@=_E-VZHgfSKg4W0(aB4g_Qg#<c5I45Z-B@MGF4Wb_CbF4(#Ad)e0T73VAfO)XJ
/4?;ZTbWPF0?8N-&P@90EP,?=;d.\NA0ZM9AL<a_<:Hg.35_4BBO^R&DbEW;4(35
;Q,JD9FB<T2I5e-E]&,-[f&WYb1<#16>;[43OJc8:g?Jg1>(D(SWNSK-[OJK25M+
L,cLB>:&eV7Y>K,][,)YFLHDU3X6)IMDd=S97N_5,Y.>)?RQM?[A:@c-J0+eU>Va
F8UgNIYF.Y+;Y-LR5-e;eIG60.41W4FDADIZ/JBf4e-<dIB?g1M<TU1K(E0]]9@P
QKaV#TLRL#GARHO,;B8YV4=P<1,CV=E9DNM-CG4:EWCe7+OCQ^.&]0HLUNPKg7/P
A:[-LH)Ub]H4HSg5XZ<GIAP)@7J3dggV.9a)0V>P>^3JJASaDC0a;,dY46G<Qd)J
<D@S(/ZgTE24O#7I&6fUN.1TPL@WB1AJ4WBCMM6)c]HL@E)D0@8c[K[<4U#:NGZV
8C+I^;d_4RQZ@c62-=[]KHY.dX^6(UC1g&I@#1F-^>KZ/gIR]E9-2@JSRd\?<?G-
E(;5[F@NSD;SY?:WHd#,gCGBaSJZ9C\Vf\V/@9UZOM-=g<&SSZ@B)9.E+14FA,U#
AIDNeJK-RbS+UCUWX[_Lf[HIET@(9S1eFU[W<SJ1fA(VG<MNZ1M^XXM6&WD[YTFG
)a\2bWQT-SE=\1NO+QBJC_Xg;eZAKfe^.PI@TD&G-gU18Z\E>AK7P,\VBSfBU+@1
?E.2]7Z=;NN?^BHR?M[TEIOBEG\JeS85?X>d1OCMGc@0PM7F46OF+;-aG[2R^[IF
6)LeB.=[>MG\&E54@_CA/FHaLbQL#FGaF7^^U1^:b7]g,X5G@9?g^)&46@YBL.bO
eLG@ZXK;?-2VAZA&beQDVAg,WB#XReEGU7SY6ZP7;^L\.Y>;X2)fO6AKQLB9)LK[
&H3W-GgMRF[7&L98;4dVc)5B^E8B]GCR3\.WU?)F1C[e/99G0CA:?/[c>;O6HLeN
LfW^a)6EL?cAV4Z=GJW]D3@GUZN][,.TecBX,[a3TYW+]XD\8LYZI_3c,26T0f]1
(VG\,SRS48_N/-MWdJB7&YLLTe0d[7cX+\M3,\C#-]P6,Y6,AN&V^IF0K6GUf6H1
@e]9Ke@BJ/\EIf+F-V62]1BGbC2X3RY>WE27\^[WM9,I9fL;c/;FA7Oa.4,<FaAJ
cRR1W>>1eMB:V?R0L,dg(IdM41AcM6.:P^NcR=/I1.?25)cfX5@H7[X#:/HHf^#)
DEL6^KcM[OVY\+12,G(e@<abf#OQ<;FLS@+K:7&T2T?Wf-:==LY_01P+9P\0aQNF
X5a5fB3YVBPQY-dTO3dLJN+GVIc?U/AUW6[W6+YVY80=Z8>?cYT8U8]I4F]9L5Q&
)[66JQ],D=2]<155VdS>#.e,FOabS@0KSJ6,5L]>.&?YTd.QD03>7cFP3;/J7ecQ
1dMeT]^X&H_U.g-ZJYT/7<6f:#bSA^G@+aG/-,>L(WHAM.,B9fT//<J?gMO9G+e6
S\O9YA^>7a1QN?K.@S(a25@APYD)f;_9)6<&3H-Rc2C9(Z>/FHZ>>c_><=610eOJ
P>]U<dGTD3RKfG:fNd(K\dYaK\=_)>g]5(.MO1C2/(a&\+L0B#5(L.VCUQQcfTQe
fLIYI1PJX#+X)V9:c?C_,3KR<DKf5-HW:/9DUCM^0LDO9PL+?U+P?FNGaV_);\>L
7acHW?0;Y):V7A9I3f[Ufe,P5C1#c,^J.IPf/,+91NZa0\&NccBHI5,3H+b7C)HD
:GS3C?.#F1Of?fLcOQ>[BAJ43F4OQTTa&&58e.:4UB\+/H0&7fYGK_dLNA?7Y</a
-f)>+39MZ&E?+,gB9L@;:ASU3aE5X#L]J;AOe@5J4LcT&I<E]<+IBWfeTd8O#4VC
SdUOGR-I(73<b5COKZ,V[8,;f],=S8J@I1addQ,9;R(7Bd&2[TL0:Y[:c3I]-N6C
.OPCKK6SL,[##2EgZ=1JW8,fbT<7bfKPL+@HA,7Y5]\,cPVU&6<#UKJ=f2c(3X>.
YW3L?FAO_B@>:3aP=>)]((<XM^2b++[YS6M]6#HDTT2#4\=+QDe>TB=aa6XLf[dK
DT/=B.bDIV\Qg5?7VF:F#V.QP78Y7SP2@e>Ef58@]JaD\;EY=ZK4X&e<95]A.CQC
(^fRIU4AL+34f>d_J(9^@?L6NecaRSXc43aHdI3MU^Af64MCdXY8E-GDg#\CEW</
Y<XRX+7Xf\gO=(C35He&F6g/Xb[\]:DBYDG:+_+b(aR0:91bBS45Nf^,SZ8N6@/b
KB93.XS@FJ8a;E:e^Rd^6=O1N#WJg/=BGZ??d:Pb7=Y(fgcEH.AdNZQM-+(N;6U_
GU5@[,CMec:L.e]Rc@;+ZEXQ4:)_,fJaA#eRL/)UD=I=S2B5-B9DLeX>W\e4Z+Z7
[\TA_<T@ZX0,N()FFfWKIcWOSeGQU,<3f/7#39c^(L(O/N5?#3ZBN.0A//d6Z+PY
EFWW@e,)(]5^d(O^1TZ4fO&8.BQMJ9;3=33()D>(2DM3R3ba7Wg\B:5B+7MHR9^5
8,)ID?=]INc=4;V^=<YJ+QY(B,=IFA&aFFf2,;Z.(#5d/O3;U;Jg9D)3=a.5^>af
DR]5cg-1I9NNe1/3cWD/)E<b-Jc34GHO\>A#.O5C^#3+&\D==Q9EF_>?([7]3TVH
Yfb/B0e)A/HD:&AMbES9Hf\]S2b>P\dP/B=:Pd)K>4,3Z4JR5[1e6\4-T+/_6123
8]FJQK\ZVN<@+@^MU0c:E<LKg#c;1XS39.WO=KP1/J<&eZG[MJ:2MT0Pf(OX]9I4
[e#BCN=Hbc(\P\.>B[E[I,ICI?QV0\GYF6_dW[M1cM3=BZg<WO#Z2O#E#J2@7L5=
F#L=/=]0g6>aK[\LFL3G+;TgUM6-;0),J@Z+MK[,K+O\dI:8M\e,YKLf:cTc;9\W
fFbbdegX=:GaM4W@>7R>\8)@2cTC:WKD._F=)@0AJM,:?M.(G#7)7<L^5H6QZVA&
CfbLgdg3L/Sf\@IR)5X.+4)@WA)E6VSB@89QW^37>:MEU)PB/.Y4,G[[4bcaG::6
-:Y\\e6Q-1\NYN;TG\NC4BdbKY4G<a@T<6F41^UTfHF7JL;OQYA)U1<RM&EIG+ga
VWX2_I8MRMI05NUFJVSK7NSV5G;P14Q9TPAJe#11W/2GV/(S/NUXIP3OV#PZ0?VW
8\7a-K1-[/S[6=<R\078Of([=a-5<Kg#JJZG2ZdM)_b+Jb50\F:T_&Y:d<3FA[-e
X4JY+>EV:9&<PPc_ZKZgIEI/>5QX3_FeNCJ]L+N3aF]UD7cCX8)=TOZaAdKOQGMa
7B:@L:(FM/=BXE6@X+Yd.+aJCF8>WO&=XdF25O[g_7Od0<d_88)9eHa^BGE+PCIF
8RVLA\HY3KKX_d&L5RX/=DFI#/-DOf)R27UVK61;cXZV#KTZP;]eF5P\NI^baHSH
@HYa&?_e_#F0E_=XVZ2a<4X87&52b_/,QN_VYQBA/B(Wf05O&G,,&.Ye]@;cD2:>
,.V(0g_8=-L(U),<d)T=XdZe:@2G((L,5<fQ1+H-]AT)=D]0<gO_?9eWM3^G(@&>
?0a?>OE=SE:Qd3J_LA>.)3^Z3dPgOJJS/XK\6:+T,2Z-TK4R@1WJTZ-0+e4GGWAV
+\01;#1T>^2)Tb_++;V^[HD+)0X)O]]L>.9d]I1-0fP0B76H3(0??ZBbWN<5RcLT
L/[N56DaHJ]V]Y@c_3OS;C8ZGNB3AP4Bc08VET&688L^>[+@d?/AD_#Z<7DB1M@2
C-GOJM6?5IFV)Sa5=B0d6M6Tg9?#+E:P_MS:fT2=)T5)F<;c+9\;a>,)#gRB3>A@
/JVB8))F\G=HFNC4aZ8DDHUYJ928=T7LDD(Q\4C+KK/<ELf(gS;(I]/SI6N4Z>cF
?\KOCEMUD>-[G;O5eC48Ma+/O0IS89V<f9T/_4GS((OD+T<W8-bF1TD=:>49R;8>
PUUQWfRM(f99@O]ZF__aN2<-f6[TDff:TCQ1R#)>THT;MD]M97V=fL/C-ULYHU2S
82,eH73S>]M&f/RGE):1IRE<4_,D@gB6+))1L(V=L#BM/EL&DH;Q8@U/IaaKb8G^
[_L/SK9M:)Ua:B:2e:0CD0Z]<R,0_8I8N88H=/CVdYQ4[SL]:b:K?H/VT@M@B\UW
]9de1CVbNf9,(aB07P(X_f+<c&XW:eC<7Q,7.eQLa0#)+OG_<Y-TEfSMU;.U3[5J
V6.C)V70+)&KAg_W@#8c--]3H(2B2SY.LD[c>V#,:Mg-9WBg2_+c_#0YTE6Ta&N@
M@Yc;)E<Ie?O<,WfF-OWQOY<+c)J3CaW=XDEc\W7;L9;D>/UgRBOLAfeML4N-3fZ
+a+CJ+,Y>=3@Q8JBO=29eXQXNNLGJ.G,E[DE,XHDWSIFQf#<Z@DD,aK\g3.;49#H
06)f<eL&O5:A[gR+=VGbIW]5EO\]_F,O0d@73SNd9@V6-VC(<1@(9/DZdEXULgdB
McE=Y]5TcJIUcVK(]0D4Y\30+e.[&:d\dKFOLaDfY8<_e77b5?>d16.J2G#)GY=P
N[O]50^E7^\\L78KOb6V,=c&R=1DgZJV@3EBaQ\.&(/[O+][6HTYHb:60RDP1VEf
fWMSGVK^<0dFG21VAXb60I-b2609A]G6dN\]M.,P=E>::VDZCVV5NN[1QM\L5(SQ
g(GM5T?/R5ZOcY-S/PD_HI9.-+@X=NYK-]HPF]=+X:.B)>eF2DI_=ZPULEL09HCf
<9MPV<#R#H_4e<d>D+eG4cBDS2\7+SWD+O+,1KZ.\@5]gLBBKBXKQdW]NF9bVb+#
6-VEQ-XJfb[?JYTGeWYcAS8fV@982XG+61G>N9:NacN&3AM>\8E-0:dUT(?X-OVZ
R@_+]YWECf&JL\bcU15=-GC.cPN.X\,<6WTX.fMON?HB0&+YgF7(BSI10?1fbZg8
>C,L72dYKLH+N-&73^,5OEYX^W@UaK\Y0:a(W)E=W7MNDPC7\WfRI-]E,4?^9N3J
IZ?#=d?^a0]KNS+(\G0gW)C9?JIS.Z-_FLO?I&4<_<R9f;gZ4T?[2DQQGOG?4Hf0
BK_3M[@Z\6C92\(-5@W>R2/69VKTfT5>A>LIYS+W.H_(:#/4:?BZ_Db5F7]L^9f5
bWCM>:-1Y)JbP:2(3W3KL)4?4&)gJ\EU<P4IXE]DHWd[1[,CM:=.6.C1e1MGWR/<
;fN>+N2^>K]=0D2WT13:fV_aB-^G\cWW223MR+[Q6^DC#fK+MY@&V,A;YG<B;Y^2
NE/=H5V6_<>JF[OB#>8gLd-SIG4#CWAc[58F4VF[F^a)7YS<\CR+ZIX_UVTN97^O
[@^7aOGG?9MUPCPW<_]Y6S2N3X8<Bb@=4BG&7;4Y7I=cfbRf.4J6YE/,=X3@=VLL
9fYbAMZba7e^Z)>&#/bYHa=4A_c97F2aQC@J#/>MJ7\0#Ta(OCM^RN.EDBBQ1TdL
?[_Z<8PCQD<&#)4UVC>DO2&gO1HKMU\CDA8R9?F,[<3?OeF?L0&J@NPC@8[:[bb1
.7/?P&9V]IS97&7?A+P\RR_)=+ZMXVcWM7+#?@6707D8Bb<aI1g+J10D5=[<6])(
FVR^7,ND?ZV5c\?3B_W;\+8d99&1#T/6YB_?+=^-/H>L-_E#/EL,,)IA-N2N<-QE
,C5&1Y&3&EP^fR1]D)P++?VL@R::)1>^W8CW?4W:,/O4BR/[c82>BT@TQWE#?NGS
F]0N7Va&XST,Y1.98F>ec)6AFb;+>6^[7Cc#W/a1L.>6e5cR<e^XOLNQ:\eT.a,@
@5^Na<L_^1:4M38NF3L=LN>9YAU#6cH5)-Q>PV7?DQ0(#7#((F\,.A:H#TP_Y[>9
<T:Ec7<ZJfB/LD0FQZ>:W?Udd[)VdFI(JJ=DX\:P2cOOTFA9KEIQ0N]W:,^M-]1g
=;a(9E9a9be^9UWD_aN#ZA8XM_[[PI97cOW7B8^4G6(Y&B.aL8ega@3>0UdWNC_e
#;T5;]B-F)B<,W1Q26I6<,(?2aB[MeUK44bV/@54I9SZNFDPSRCF/CCS/P)>D\D0
bJTNMZ5e.:.M@Q86BK[(6M&?_9,;e=bQ?;9>+Z:Dd<?bU9a&D+HZ86c?UHAg0)9.
[10M]90V(Q1gKP0X5.O]M+AR\?_OUGVG(;(7-0O+>0U;1BENg8F;\6,@cD-W2CVb
(d(6OO1HADA_\/1\Xf3UeI#f-g4IV_2Mc868g([eO?;b6Y6B1ME4<GH1&Gc#PbaJ
#-8gdeI;P8D:G<;VA)8I^#/7E:JY=I@](+T[e)=J#+>f_8FHd(UD1((5J;04P_WQ
BfcV:#;]UK1c#?<UY0M6J8H-4U#90^B_]@,,]b;;)fO^TGRGZe-7X\6<S;:]G?=C
NcE(6bdb#1?G_OQ.@>Hf4(7AA[a3X<:,HaRGO7WYXSNH/IW_D_6McKS<H[H;d?Zb
;5.4_/)N-,>#ESXJ\L[;f9\:C2;g__,)>_RgF8_@Q\^D/UQN0E_1I)8PdR#RFR)e
/&ZK33D0:GX2EE:g/acTK;8/1DAaC@adQ;JUUECdaX]U\Z5_=/M,4JZO)4JFO)P6
GbTYYX81fcB6Jg.?KZcC:WP/8C6(78EfFQ0TRd4_BHf1,8@2<41D0D#\bAF]DWR,
c<N=)Dc_(EP?)1c#K2&COF(c3SLZU<2Be&DZd@;Q4.a>8V_>8_0b]1S&6JW<O-A^
eL/VZ@&JL-15@[8Q7[I6I7a9>)1;c>9=Z?4XY1T#/X>=P<+K0.=)A&.=H\#3gc2B
0R84I-WP77g]b,MASVbT1Zd.>N/95)5:1:Jf_(b-SYI&b<PR)H7Q721U3J[_2>>_
A-O,V&^LXBBV&ZE5OM?42-TEb?@W5fLU.C(CE]C;JZ3T(V,B\84T.+4B-&#F#A^Q
85D]Q,:7aPBZT-bW?\U-D9/2_#MJM4[X?V,f&#ED^WAI?B)H?V\2DD^\fKQ^SBN4
U0A3\F?Oc[2HS_dI_YGC+4.)G0M:9RE,/GU?\7U&+XD2.eg>Z+90D<GJ(E3LG1eS
CdaKR)46g)Afe8cUgZ(b/X^,3Xdc0IMJD^[\ZQ/F+7H^=/BD[HaY\F0:d/CVQCK8
YYNL#:9d#a4AP7?]&RQYJ&^acZNI4?Q(W2GE[LBVN/Mc#X0a1)31@W=X]+c1&@If
;R,#P^&c2TP5JJLMN9DSe_>_26MYa_2IGf;0gc]D35DL5#AgX8Adbeb#/Ta_:c3F
K/9UdKP;cS?57;-;8<I2BZK?X>5J995&#R,XT>RIHRU9ESBH?Q^75]K9VgXdgIcY
W+2KW\CG_8<IP7Z2)bB<Wc>2CZcBX@Z#NIKC0GNbP@<^=;JZ(T.J&.20,[V@0O3V
-K,#BN/?J?5?NZ2&/<T5^gc#V(6@TKPSWQKZ,N[a<X&>9UV<_Yf2fO7b9K=dc3]L
77W0ZWCgMJ#Hb[AQ<[/78bA8/6O4NLD10C#[)f3[I=PB:(OP7A&R+gVD^ML4-HCf
CD+/#,+,?PXD.0QIQI)6BfU[33EZR#DS>H#-.&,8eFI@=?YHO\(d(YRG[UZ>]/DW
T^gf-<[Q2TJcJYW4C+b<Xc.0J=;f=dVc/O@2O-L2PAC>C-0&6DgY4&ecT.S?)cIe
>^3M[We1O6>GNTJ\KPQFV#S#4+V?[=U8e)Y3F4.gM1cA@,?R&W6SO[(T3MTMT\2A
7Z-A33?;(XYZJ-FQF)dCTSJE-B994a2_Ze^D#A;NDD?0Sb56EZDNgP1H7Sa>YVcP
WNeLUg=(dN-:1dK,&9K+?=F:6NcVVUYP#&B#J+K+LY<]fRLITd+fM._#X2Z9MZ&P
D-dV?H[:2VNT-I+]C3NbRST-c6^b5g5A7Q\X,AX&\C?fIUR;8U)b:A#.WBBT6SW1
Pg^ccXeeZ.&P&]gSN;5[4LOcG/71@1I4[]?HN/aT?<UO]9WYY3Y+H=O4)V&Y>JF3
/V^7gVFG(UEaWBe):]EI9B8]))]=:[=RH<KLFPXTWYUfS<bNA)R)eC\9dKUfO9E[
[HE+G8O]bdc)9/T?Xa_<Pd.CND7^(-7O8(X==2L4X^AW+B->-+902b+S,\:6VUfS
VLP@Q]@0^XX-J#Pd9ASMYUZ(@#&W^,(O[J34V)53<cNQ-)-CR3Df(>9?&4bJX@CN
DJB_#H=<4^ST>B[=G&VTLJJAd<:Hb:W0,(/)CRFHcC;EVZ.0/b17MO,2:_cOEJ5Y
3<8VJVXC<Q67c;20c_4V<c^DQX2Z>O<?Ja^eFGKIe/gG\MZC,T#g[/<Q)9UW(d<2
=7T0.,T6_/@Db9/+@Kd:^^_fC=5A_.@&?9(X:O=TW(:M/>d)A_#aZ#>+B7_aHE1T
/4OKQeAX>XS18f6KQ2DB)=#e&LHXBJ9ACcg=1&4),2(UJgT5;Z@<gEA9#2&U_B6>
>Q06=(BAfKe<=>9-.9^Re_;CM9+OMG1)6N0/5)A#gC)(#aNQ&)L#;(JX3;<R?9LG
9#(TSI+.B[PVVf#f98PdIFF_;<E.Je+ZRS@4[d50TMUYUc?@+TV)>BEEP7)8ddHW
8b3_dO:#)7:L6Z5U:YP:;Z973J9,&:H.F;NO;W@?3=3J2SDLES2Nf<<I1M]1DKdf
,YAY+_X[9J^SJ^M>d7P]XGdRJ.gPFbTacQ8ga3S\?@O]+D.4#]H/XLSH9V,B\5a8
<&YHG<bML<d>X9>.BT>e@e0Z#)5A[Ubf4\_)X^eY6KfP8SIGCe>T9ZX&&4;YV5?B
4XGdW&G.M3TeD87N;]/]ZREJ]V[BFYM^YOcBfEf3cT61D_FA-SG;Ug3/S8,T[;B9
13UUX:19dHR]BE+9R#;0dVGPI?L<)//B-?)>/KFFH-MU.W[bDIUU7;a0)(,d=>ge
Q+0N.Y[8fNdP@,G-MQLOWV#1cKU<S,e#[BT3e=2R(5E/?Ea<&U9PJYKIOGSHgC8J
/@5:/HUE5O/_Y8HQRYdNb>C]H/dS\Q5bKa;#2CB/QA8O\\@12(A)>P+Ud)J(<B_0
OEW-F7UJU/;\MRPPHfD\U8e7EF(^A=1+\J>N59.1TEEV.#LE,5eL2<g.AcI)1;Q&
-PZc9^.?L^cRd70:9;Sd)8L<0S6BIdLa3Mc-1?9c^V3fH^,FXPfg1MFPABc/PZEK
JKBI-EbADc1:O^2N4J(S]@g2ZV^gJ)SAKD6\;e&f@_g<g#6T?aU@^8?9f)RWg4&?
KU;@SPa+CaALN,?7Y4AY=RVC_cg9Kc8KI#FF3HO97A7S2VJ6]34._=^AP#D3bTG5
,83H:W5BDIU59daR4N4Q&gIf6E.HGTTcXDR?61]_QZb4W_55CRVA/:+<3AB21Ye-
Y+[&faHD=(V<B]?=HTIT2IUF9SJGZ(<:,@S7AM6HGK6DXWRH<W:0c26]aO,^U9]O
SgM^O3Q=;IVIFf[VJJKWI&X.a96+JB3[g<=NNJ#VegQ6JFIQ9MSU_SR^ePf[?UFB
cKCP()2.+5OA)f7;;+O#gTZ:^/M8=PNZ_N8LZTNd6gFHDM2N]D<a8BNf/(&:a6=<
<JaR^5-EH;#Qa^0O_#]a6dPdD-Db(Mb+bL]U&8-^U<I&E&?f59<\c3ITScJYTM3a
0:[FY47J,\3?ULD90)^eE:d3;4XRYPU5RB9DP5V)4Z6>[\=\Xd0J[R1KeT>,>A/K
fbVR1#6.:>V4;C9_#Qgg^_,deN#J8;0K?fAf=WQXLb##+QH&V,Ib1T^CW_6@C>VJ
130E2254g6?U@Oa^@Xc5O#cgL-1F5,&OVJX_1_6^W&<==\\4O6[-EOad.gg=8DFe
c1\Gc>U4F)^[-V7@_@P?JWBgN>X&Z8U^93INGGQYBgOYJ,RJ.]GMJ/ec&NZNB70P
Uc+<)Z(8^X36MW;=d5f9b=M&LA.6P5U8g>f_W^CNg(1P3.D7D1.@&B:A(TE-[:U<
5&9PQ>4Z/_(b8KM)^CJK5FA2aSLKJ:=_WH_;:^CG]]fD+[<_4YQ06UTBBF[8_OZI
3b_FW7CdZ7Q(D<O4Z([_9Cb:\-9f9,]Z?ZdL-)XfNRQB5-K&)f<&.9?X#P?:BE09
1S@HUbQZVaD9ec^LCgF,X2F/+b+ZUK[>//<9a>LQbP#ATdVgPT4@/K6PDC7gB];N
)<8RN(Gf(EIH.NIK\&F=HFNG+Z<bG_(DZ)<WF4K5H-f_U]Sb5)BAeC:T_GS5_-FW
0-CD\7_bOO@/:TVV_ZO\Xa82JVX+V/9XH]VFC;JI7T:\@:0GK<P>FCBV-C8e4/..
I&;,WP#K,]dc2\[S9-82OcWL3,U;9Gcd3LD9[/WA]FKgS^.AO&Y#_-L3G)J+eb<+
T>NVIB/T#)#4Cb?(-_:#/)4R=F1SR:)PLC2=QKNXK&GdG.DR^P,HHK[Q8e_&E^96
Fd60;RNS[HVd^7)<_He]?Jf-0IP=^]2LfV4C1KURK#^R/4@J9ZW/D>B>LITV9aG#
?-9aY@KgBI\cVEJafU9:8M465gB&eI&[dC1UWQd6+D6_1RQ?D49?&5#)IK=W^@93
&ROd;\;9VBJ>>7G:#Xec.b;\I/8e>\:^:TE@Z;.d,XT/,[PGHIUO],-N(HXb]8Od
3IPdCVY+.F8ZP?_eBH();[M#AO:<V19CB<6<U&GBAQg2KXd=M+U+&?:=DT89=Z<U
\-=\7#FZ+;CAgYf>1&@+877Y[GBYJ6f+6gMO6W,]F3^Lg[@3)Z/@0:V:W3D(+=<[
.La6eg]85BIV71SK>&[4RfA1+@Y&E5S/.>RE=9g;aLN5TK45Y+9;<V5@e,Jd?AL4
#,)9R_;H]+bJ\[VQUUF;LG46[EP8&V/_5;b#:_W5GU2L:6&0C.@#a&^_P?0Af<(M
#W)eaTUGd=U5[9Y&AX6@3;;&AJ]A-];;9[9&@POJX.Pf4:129C4RE7VEeG=]/3KK
LHNVN;e),bLX9#V1]2#5S]3-4<=55X>OA;[?YM#gQWE\5_BcTXJNBacLc3ZQ+8RR
;<9MF4C&0\@4bU9K5T/f[BR):QY31#gLXX&WXJ)>)^MGe-L,dE+b-CB&dge9)X2\
DdgXK@e:I+^&12Bf97Z[0aA,[_SOBP.#&>L+fXa_W(g.YD1\1bZ\b-J<e@T8\dF_
OfKH.WVDGMSIEg70X2\.:S^L#R[I-427?X6<9BTBZ)WPEP9O,KJBJ8JC)f:?S.S=
A)DV]Aec_:1,&Z?gS2TX==.Ve1)cT0=P2RZV>M7?-C[TE^=]KdH6NXO/-YDgEN1G
[D,<8eb2DEQSRF^:Y348fD:&PXb=2BW)f<UUK&_:A[79GF6@8&F=KV_N\Ydfd6]Y
JPOWX][0EgZBEJAd.&A)/>f4,,#Hf9SH.Q0/eP#=d/[c_#9]aa>UJg,:8H&AORT6
L#6<)6@EKdfX3#8/QJ-F=/0fD[SN3+AVEd?<7gVfBfLbc29YRVNceT<>P24:?KC9
\>7+<MM#ALNR??Keabe^^^I5#)HU?[PNN3KOM1L#BP5JJ8S[d9=?beC3CLO<)YMf
3(-g0(d-(deGedNbIW<#&VNY7/=QX\.+7L5O52T8VZfd&(M&/A0EIbLFQ4&&:1,V
Y<@#)3WBLfH76?&LKbbEEbQ=[K/D>cK:QMU/P&\)[#>H^-Mc#K?QBSM,1V14)b-E
NcK1fg:cH5g/B83JM,K3C?f#[LW_2;&>(e4KE0Mf.DZ/2C7e;WERbPeYGF;OGW#_
fNe0>/;N#]52=a-eI3Wg.c_[_Y[A&XHZR;@Lg6JP:b7Xa9B&:FTTW51OV\:QV)G]
+H9/S])(4K&4KfGIS]LPNb\M8QH5]@P<-fV[#f_YD?_;R-Y<=c]W\C[6f,BI0680
9+R(DA5)R4C:)+dDE6=^T7F3FLIgVRB\eMUON0]cd+?EgU#X/g@L](K/#;=+AFB-
#ZbJ3BZIF7b<#RQ62,<KQXZ1DGUZ:G+U/.#Bgg<V#IUHEg25MHY1DG08QW@],WKA
,YMQQWDaY/+QF<JeHcQ+?_CUd#MJ,/8a#J^:@7L3dK_Z&dgd33e&&bG9<OYY<eZ#
Y/+4C(b#@0:e+)JZ5JXQ;?29gM-IFgKQ?Q;59LV/c&?RCV?^3=]JMOad^+<O7O=Z
,F&M(Gb[0eT&2[\:FOHV_.SN2U(1HU@Jb;e8AGXE;,6GcFGf?GG2+Gg+U6Tf?RE;
#EH7D/LDT5FTScKJGJUB\9>UHYM]1T?[G^.+P=X06</Tf/G/DD+T[(<WO6]H97M1
bE5Q7<OMDdEI4WXTCT?]f[]^:,GaA;7gDQ90-E4JC=7C6OSV5HP)OUW59=YB#^8A
,/:OcX(Y,:+e\YRDCUZ6NfSJc7BZf#eM>dH(\eG-2W#_NN\U7UgC?b+\8W1dbcW>
fA_@Vg)V>S<#C8PQKJ>U+TF^[:WeE0=WAPD,LaV:&4(W/PTNNeWS#Q8)X-CKR]F(
/O,2Z=aE<XPRJXLe-0aUJ@]>Ldd.A.aX0R3>#G&:fXIRff>?9G9YR-WAV/g,>R_E
M#BdB5MEX#21BS(+6dN3VGT(,PgR#U8,P;6GT,VTII?,3W_,e318YF]E8I++N+YO
#:G&/#TZV<#aGRAb8G&?-5H?g95A3eF:+)C>=e]]9X0<>B^T?/,g,DDcHGe0:/E8
\+b=dTNafVRJ0/d>J)NQ/]7A4FY1.GaCWV/Z1O=?+1C?[FM)M[MQ?,X.aMgC<XKU
G(eZI,CVf<2K&4.XK<bT9Q5[D:EDc>VZ\c5PR6<(6V/<DN[0G_CT?[_#8AAXc4af
L9dBT^H8=@Se^2gGF=Je2XZRK>2bG,H7@cM)GG@aLJ]>ef8:bTXVK.V[MfKL99_E
A:A5^B@e+\@gN_,2Q8/:ILD9IV3EL0HZBWTg/.2H0;Q?\VdX^G:HbY&LU[A0KG9&
FE<d1/L,4H0,10^Q-U::@@90fG4CU-CRgT/.HY<d2^T3VW[S<\6)VbL?J>gf=bAV
Ed0[UXB=G;/>\G@6X\?P@#588:L:IE4WY#O/Xb2bKA\/47a1CMM5&8TW](0IY2PL
(7f6=0aY.,f:11\GeIHDc7CK:0F21F(L_GbeRYOMDVEaZXTfW&Y80(DDF2gdfM>U
,>aIR.;?JY;:4+V9EW,KcD\5XI]+a0fgfAJ-\KRO7/3aDccSc;e)7ZW:JNaOYc-#
97Va6fKd#9,QeMBT:cN6<2UA?:D9Ja/;&fdC(J72;1>E&.?UM-=Q73/WU[TB(3JE
c7H2+4Y,,b(f#J;_L7#c-,52T7<,B?aJ#8YTO/]I6H]P:eN2K/[,:<a)KLM?R9#^
A3.ZCf:W5&>+&(7PX[\W646O8K\FT@<Q4HE]58-R=GBV?>[bU7.2P+JY[<?&_GP,
U&De7X)SAC\F<_CT>aX<BGJX5XP98:V6+^8>-VG<I(]#2ac1>DQe[9U8KdP+]C?<
SdGZ_\aJ])C_ECZ&L^)If7@^f3cb6&8XMX(aDFHGF:1&Ne6RT9HT++/[PROaV5a:
@4a.<^T2.;C>6?3V+@5EP-gRXCd((]?P3K;\&R/aM>J[aD1WS)X_&5eM_=DYgV<O
VVHa1-\NbEAK@FIaI)Q@54)7SY\MZ7_.R3ZE3;d@_W#[BE0NDT8B1Td[/fJY^X&4
RUV/3-(O;-Wa1(3Mb#Td&MP:ZI>VPFa+;444JS)SKOU-B4Q[\]_93gc+BSG\0,c\
fE/(]>EEY#E-)VaNGd7P#S;Sb@CM;H).&D^V)_g;ZJR<@aQe.Q0V^f)O66_.AINW
8ZXLZWN[D75;TgAW562&/CM;dJMGKE988TggOV&F9JC>g[EAeE9Y=+H<E,5L5X@8
bK#I-_/]A=Ab=0<P-ME.<W@320aC)ZUF@FeTY2\TdDUTVO^_bD7[b1AY18W8F50a
5>:BZACaN)cVfe2&)\ad:R9R96AHN?S])KF/6[-<ZM5We:Z13OK9K7<4M][XL/Mf
Xc0BCOQDb8.^?,g1D)GSN,fI<LDHPR^PR#B/O1_-KAH=,/W=fe:/,)5dCO>9^1-Y
A&b6,)@VG5b4/6RQKM>1Y-7:0W.GVVG3L<9b=MMEB,@3QAVLA[3:?LZaIM]IR@J[
\E5):2?DE6=P;\;6+/Cg]?f_-W</EP,JZS\L?gNTP#C8ECLJ2Q^^b^P:1E70,Dca
;4^^VdM.HDQ6GPAMR5)+ED/N,X>AG/HW_EMXAcgZc#CKUa/b0LNW(\0,0YFP(,6F
>Qa0(KP_Je2T\PW_fTY<7ELL<T8U^@02;+bB5>[M24KFEBcbGKS-F)O9&,ea_dBc
3H&L73QGT98&V(]]@;AT^X\EDN4V-&.B&-FC+2HX?c?ZJ2/Ge2.[Q);CPNe^fVQX
<>G4Y-af>2R#D>QA;.?)g\>D7V],)c6ab1C9?5V=>Q-]XZEF>dH4R#&<X_:Zfe[K
gbS(8VTPKXF3:eaA-+M0>JU6MV9M7MQf9cU=,)MgU0X0/Z4@)3;?9]E-V5^HGVag
d<?_a5FU5ZMHTNL@C>T69#/U+gg4#23&YYL-:GN6:&c=GeP=7MSg)bF=:c#^]#P[
58gVZ?N<U+&K[J3R#/.2(PYaP5b]-7WEIE./USSH1F=.W<,S3&W,G^:f]bY?;Cca
0&X#g0f831?PSPS7YX5aNFd3X8N<K:bC;N81B53Te8A).=9HIE\7L_A\A3fA;0eg
6_JI1^<]K2aO_T?ZR&)UC)FD(>aBN/LS4SE>fI+5SSSP<8g>M6&_@CR1HA;3T@Z[
KQJG]AA[+[bSY.K,\dGL\FGEN4&BFX?0\cO-M#COR5-NS:@@O/A1bZ64f3)e#3R.
.XeG4Q[G>4^d2W-#da?X?W.V8U81;+Zca8#2bX=:fLg)KP=VDNL,@QN=2)#HA(?8
Z>:4bW)+FgT]OUNH84L^15B_OSaPM<+4&3OBO-OF=6aK\?N_G5W2J6PIVX3)?Y5S
d8ZQ+Q1^_JDBF?RUENae@Z(fQ2PF.OG77A1E.Pg6KYe9C.\=;&0aIbM5_=.?;<X@
,&HH-X(eS7FCFU01a=PCf-CXC;@,=XE5X^W95F;a&934cdZ?Y[]T:D]^)a?/=[Ug
O#XYY=+UVfS.fc6V75E.f:f+B8T@f/89#J,@X8a8adU(WPMP?UE&?,^#eAH/58Rd
Y<?OQ+(:@OZ=PU+_fK0[6VHJPZ[(^f7_6&[^T\_@WD?M&[<6.BI[VYW?.6;T2RR;
3,cZ0QP2CN]H9O.(2B1\f9BJL7Q(BL7L;W3CC4AR@b>UcJdV+1A:H0[_R9fE295C
12?>5]/M+/=?c/1^)LG8:J.\;V]EaSXUGH[AQ>:&G.dTdQIJ-=,/LN:37,Rb<D>.
L]>SU,_f?8SR81-78<STSB+BY[EYdc)Q0B&-E<8YYZ\3c#+R]&&40];WO/b#2&<P
L)d&faZ640\f@_dJa5bB\=B8fe09,&dbS4G=-G>Yf7I?OIWfEKa=.DbYW3]1,<R-
GH)2#b2M5Q=7d?HT4P]Ug2Q56OGUN&]Pg?&VM(UI_7M9;d,;U+g?B9W-.-\gf/)&
?L?d75LD81=Q7ccX8[>(&/16#\@-H4CDXJ>JS)7T/ER6;2UG<<I2<3RN9:(#\[C9
)FTM5U4U5+LgRJ&Nc8>X1-3<1QW)YRFVT0>3]&dMC-A[+H??<7DFPESJXG[]BJe_
#HT\U+cLG325B2e_d5MAZZ87):ba>DV#2fX5B6XXfDT)aR_dLe+IePg#<feU8,D.
c(K3.@.)a,?2^7H,-BJbEMGf8[V?Y;WMHOBN.YUeD+Kg5cgf\b^(\<#KbL:Y>UJd
/R9CI0I+#QI=.\c82JCX4ad91dagL&U-]AGRHP1X[#FgHUMYaX@#]:U(R@Q@F5Mb
]F6e5LN2E6FaTR#,M@YF-T:)V\KKTAUKWSJ2HeK\@,]O]JLZa0:OM]bROYT#@M1c
GEQD:6YW?.E>RH:/IOKa19KWI^[C;+362A85:A1eZGFL0HRNgf-eTLfL1>)Y+GRT
.c<]ZCc,Y>a)+S4)Q/e[OA2C#^4DFQ)D782J#QJ9;dR^6U87(6EP1a;#B4E_0fZ>
2S<aSBg5D=31P?f>PN&7KUI;Lb>8MbS,DO1LHOfFR1PR(g=#]+3_7Cf7?2)d>(P/
_2d-;S.;/4_dEb7FO1_W4<9ITTS3-;=(82d<c(>I^Pc:Kf-.SKBcDP+SBVQ.f7V7
#TN/(_e]QU^QbO4e@f&M(::FP?#8<aPFXEV92Cb)Y46d#8MdI6e[J5]3[DB,O:NZ
8c0@_(ANFZ_O,5NC8gI(K_FCQVcJ2g5P7ZcQdOUY(X8U_>cFdYLCDTU]O(LEXe_#
O5:2@V#?-W_\2GA/X6X#+FT>;_J9&/[>71?2HZQ2L;1J+#-3?09&13_V[P(45IXe
.0G8e:FM0KLH>:8bNWFb2DNf\;_+3Ca0S@47VZB,HbW?XSA\.J-Pa65EB15C,eLY
5I<a^eKK_VdP&a3G>1DBO<,HSEH<^SSJb8GTF)OSS7VD+:6=GI);b9&?O0K,I9[#
;.SM<MX3T&O<eQK.FJ8bVd\F&6O^5O:(S#=Y,+A3()U#IMM>1+C^0U.H:2K1<NU@
d_>ABD:44Pf]->Y=bcCAMNS+(LHFFA;ULcMSIf5d6^KCePP/Z4b.<T^P+a@?]VHT
X8MB7G11.D^fdY/MfHUga7G?TfD>:^BS9[@.P<):=V>_(#DDSXJL[DA@IKeL8eFJ
/JCcWUc5\eS4[XcNOeS1Y(&2OUeHP#:P-Cd_0>&HDQEB3#&03NJH_1FG_?LSS&?G
+Y53K@]LV.)X[-0_HKD7:46bVeC3b@B##Ka,6PAJaQ=FA[U;&/?O7_+([JMF=[VJ
SW@aL.@NU1D<D\,4\#cH\[1HCT5YaKPL6HMWRO(JB_)1>V)/,1#Lf&^O@K?+f=SF
,R:b-97+JaMD8B<+F[7R^L[O<EXY(.c)0#eUT-6YbI-17P1U>Lb\GUHF)&JTCRLB
COY-STX2LKKdY,F+X,Z(e6Rd2T+3T@J[)e63EfN-G4gZ./C8YNG<2<M4LK>PN1+^
XZG#RC6bX=<0CDgQ[TYU6<VMAg]_,][IE6g1&7D[PLXaJ01?2=18^cZVTPga#H0G
S32C77DO/5&f?>?<HJG=1,aS69;1A<BNOaDJ#G8+K^&Kc7cKf?FI-^9aK<0.9_@9
CRAaZbTO0YV&BgUJLMO&,eF;@4f#\&&75LHa=1aBdf6D=M,6WT2GJ15J9<<0Q)/7
[)5OI_f]S-E;A,8,^G/=T^QZe0YL+7GA[Y5<5gXd<Q8JF_Y@3\Ta9g(&Hc=6\e?3
?>TNDO2B<D,)594^gY)Iea6bRY?L+ZLI43MdXO\?.Q#gG1W]U_LR#&C-X.F-S,HC
a(T^4CEcSG&Z\c_4IPYcS8R54C-#BSCFL:I=-=9,TJgKV\?/TZIaG6)[GXTN@^53
VIL5XRVcI[Zc5QYHHZ8Ge@03BcE+8O&b)^?MP4B4e];4EB7?/,7gb0]J4#<#XgCT
,VD#\[LME#+O=QQ+4I3^Lc_f;VNV9-070LR,]aMFbP\/a;Og=)\/F(cEOT^,.OWC
25Z7^A<bS:fMO6@3Y,8L#R@?Z:J5cF;:f;98XUVN5]<5d20#UAXY5a7.C5KQ5K-[
SR#?#4AQ(&8[eL.+SX<)&a[=>E=NZAVP_7[^=.LfS]331MB<9PH,YU.OP3AN0I\F
8EJ6O-^/#fYHE;dTQg3V-@+WEC@OcM5G;b9J2@-#2QZ\F\_O5/8=C0^M#QKZ14Of
@S<MfTFAH6K@R3#.,g]1UE4Ue>&5TZBEFD_.IT,^LSVSY,H-Y:]&f\cT;B<?0fQ+
U_Y1+?E>H.J(E-)[+>R<c0eZUQ+FW)cdS<dg1(>Zc4L\J#6W0F(-7LKL]=]ZUP2B
AIQ@a@>]L0b,.1QdFA^d-YaO6GG8O]LEBG_4gO16645ODSZ8/8]&ESQ=J]W_RBgR
g5MOF.CAVd;)2d727QX/Y1D/T\1?YA/4-Y?TC>CRDQ_?0:H;VZ/2e1KPL13c<:f]
\g5W9PK^,7I_X-?M<_7^gKYb-b\S<NPf\WUT(/44;]2GYIN><<^UI8OY6aNfG,S<
>04/G2bS1AffE(]H<,?Ne<MW[Z;(4eN]X5?EP7K:\@>Z5CZcYY:_]3MfCR\[fH=^
XT,dLTee?++-]W]&1[KbfQA@e/:_^/a.N?5NJ=A.6@)#0/d(#C;FJ+U<AH#HD+IN
;:&_eY;8&G328A8#+@UW,(JDKM\142J(,g.C5JaVV2&UI\:bJ0BH]4b]a8(+N(Zc
TH0,(--H_E[_TDNJWA;T8]0(<AQP[<7f7#+CD+I8NT/3)2F1I;U>5PdMC;N@(@GG
&IZ7d[03#19JM(:&\,</_HDO;>3d@5Ec//bgAd6+C6GG^dY3JZNbB#&XTC(gebR,
5H9Kc]=fWR.QX@I),3L]ER\RD<ADg80+(HQdKdIKcHRGZdS7P54R6J7Uc]F:ZSJR
B=/-SE2@eA;c-=JW0G/;),+O5VQ;4ATK:J&6KBX.RA/#cc\L+A8Z,DI/YW6,SW04
Y#UP=7RR=ANcU[cTaNdU5b],0=M.61USEc8-cdWBG.5,G+@ERL)E7OA,a;,#WJeH
WJE[9gcQXZ2(X]XP(/W:Kdc9d4)4^+HeQ3b1VV5Z1JREXGI_D]76+T.dIc,;Lgfb
Q7R/-I#-cCd^O;XT\Q,T@IN=eb;U8\g8eVBZZJ:D;)D(W&Oc7?=B36_#0MN+Q+FA
M)PVHbD+d,#c09&QC-F?DCE/]g^N6^0/U[)a+EcH)4@8CY=ZTM(Q/TGf(35H1f?G
UZ\>a;T#-?_;cd+V1A^F3.Ed=YT++O#Z[P>g[7dAB2?KTJ<Ff6gIBb9DNT5?M45D
X8Xd?DL2_gI]H_>><C-AcfNC]MBDKX_CCM0B6f;MI(d[?U\>,LJ@3LRb]NB_4A>e
IYPZBa0(#SbJ/d:+D[\--Z0_P4a<?@--J#Ig7Cf^@;NHJcD9O\?0)XB^J7,6<P]0
,9;^:CSMXc+Z>LIXfM7)YGX9PALC>GYEQ8(97H6<S57X&#+EH7D(\1@BbXH4]S;(
dP/bC)82a8AO3Y(Y?W.d7BcQ.00JO.SI/_eK#-EGgSNGDO\7#,XRTL(,3E5FM)DE
0[S]M4)FF07TD4[?5Dd:<B66UQWL[7?U;V?W9<Y)+;]WUO@ANcFF1Ra^eS)g;8<1
?^f6C/GXTRF)+R\Y1+a&_2?Hg96V8Z+HgGA:<XE.[A,[GXMDcfT)J][>^\_5>]QO
9]R=3WD4GD\Hd5E4^>+0._gB/];G<8C?IBYae=/^CKMPBAA(]I>>daT).]LM1gQ&
]_2[d29g[G909FZa3D\B:JZAUfdddY39#-Yb.R.D]bDK;;;LZG#d&X41)2#V,I=>
V;b&X(:F8^#UTFWdR,23W:[\aKa3U8dIOaB-YW];9;1c#Y/U7C=GgKZ;&a.;JW?b
_FK)2^6@@WYI3Q6c+W.YZHe(b&77,3-&8;ZLAOFZT@3D/bI1e-B<=Qe>+O]K:ZVV
eC5;a1+Q^1-LMH5-faWYS2IH1/O)ba6<b\Z)1/?e5VC4Zd@#PgJ&g&8S)5@]c=e_
N_bZ=5@:X\PWJE/Y[ff11R>V#V1A)D/cg62YXagOdT.NUa6]3D3TPR\UGI&]>I+M
SQZ.f+:,U)BZUHSZ2X25J##>>4H\^KJ@9c>Ge\9V1cTa7-XLD)VT2OV<;.U^N+gV
+bS44f]bM>c<Y5O&2GC<c#(>I;+@bK:-Sg8.(5=;7JW^=fK<9LW>>XUA\\b?LA&1
^UYgc3;EV<P6T18,Q0UO+SE.7L,=@TFaWND]&7YC[,^fY3__B)]NJY3Y0;c2A4W@
f.U-/f_2eU+DgLDg\N_9bNW^.]#)OJe\1\@.R#MV4DcVDOfUeX55,1=97&H-LF#?
4L3\g82+ZNBR\e:.2PNM(c4R^#/8,>g4<aa._-gZ68&9&?ES1(PGFN4;1T?Rd?OF
UbWVBg2VBD0GZ,S.2dcLcgY[cVfW+#F0Uc/H4L;N5Kd<^dSFZ:F1@aGccTZa+)4^
F,QF+e<HT0<<_45A4eOT7:F3b]:d4fG0b:&/9K1d0P7D<J1ec4)R-XF;LIMfG>aZ
40P02&4aY3RM>>VS?UcNcb@cLQ3\8XNH[9ZGMJPCP\#NcbU1bQ9c9;IGYM3]X6BE
O@)GCb697]=(:SG&=SQT:))::3GML]?H:<:_aUd9T@PZ^,.&Y3C\-U@:T\KaKQBK
,2g)@-43.1[>]=Y0@>5O9#M04H]GCR3NMaG]c/:=:Y8TK\KKS-N4UD#f7-dL[<Zf
-KFb5Z-D781>O^J4E4IddL-W[C(V/L0aZZ&aV0CL;X[+G3JZ8,U[M-:70_]ZeIAZ
88S5dX(T#/aVa9[K=2Dg6#fL8A.CX@ZK4IVS9.H[g^(=KDW;QW&-,g5]+LF(H;W.
cF4RSP@+=.D)>>fUI4H)ZdbIe0^V\UOYLQ.-;&Hc&MeL@GK+E[NAQggD71B@E_Jb
^)/IcJf+&,&@SK2#\BEYYCF8=f2UO]DbcVKYY?I,GZ#a?0VKV#9[Y(7[O<VKQG52
8^MUUSd.?S?1=X,S^ZX(NVSQJ-37OBI=X1QC2OIXKQ4M;.[C\ZB^:XE5QSQ]UFId
(0a/3Q^THcB=R0VB;K1@(AVO76B&GQ:6RFXVK8AYf<.^G2_EMM_8QD=]cP+@=TFU
&H6.)BT]U4KKF.eWQ;,S#Ae^>UV=)&MK>U0[=23bBG0[O]240(A\SN5_69)gTQ&X
_PO/Z:]?/+;g./MLcO>QGVH[5+O8PcJ^V>EMS;W7>aBaG/-K2fL/80^T.4\==Y6<
39]?cdCTC<58RZ8A27-S9<,6)aJ^O=2Ofb+/W&?H(T-A@N[6B,X61.c.W>7=]8D3
(gX:dHg=</+-A=,R2Q]FL420,Rb9W()>)U_.Q[+4Q,V6F\+F87^g18.Dc^0[EP.T
9/)+\MX0bP:>Q-S+fH>[NV?XF+&2#?WZDeXHV?Vbe+R-5W?[/413[,1f:-K\<7E=
,Ub,1c;gc#Zb:55:M(;8U(+Vd5T3G8C:208IUTF;d4E8S&V+^?#E=8575[N],ad)
NQX.c1A=L8Q2fWS_?6e5a<3eFeH)3\^fRa](Ce5>:,8d7SH>YNGbN0;33D1H_f/I
5gd+P<1F0fH-c+L&#3g8RM_H5QGd?4#<?<+U=VOT#H-YZYfW6SgAFNGfIP(U0<63
bB&L3Y91/1UP:&:eRN-#&)DES3f^(d6)SYRD1#\=dC95L/Y\CX6KE=:O&Qf_VCP9
M@H1)JZaf<B-]KYX+9G>D8ecYbKQ14YWXgUWCbTD8^WL^FSFNUI&FIWf?41H#aTf
RN_@25)JOB:Zg_J9W((@J\4K)3O5I[9E<cEJV6T66+bJT.,TY@)>F#-@&GHKGVX,
:1+SA;-4TS:][^X]gf5&QXXX2PSO>Q3a@L8,G@@ND.<>S3UgR9<7B07O.:I?Z9b@
OQg5S5eYKF/e]XH5B/U_c1cEWe7(\,=.[cK)=;VeRd3PQFE<-L\=IM8)VeCSJ4:C
,Ka76;H[(U(Z2(;9QV9RR_&dVd@bZ;S,Rf\b6083[B+@7]@Z#aBF(@T+M7OF8E@(
H_.CIGRUX&P?A&:[Odb57YOZ(_EOgb(>9>0:I?6(9\WO7?676(g_)Uc3CDW3O(;X
1Q=><#0^.XV03L?aPT]7T@0+IdR\XgZ:U,7Q0f]H]#Raa]EAM)UD]WP\NN2RC]aS
)cZ#&\VcIXO8g;EJT2g@+,KgZ>VbNe?MT1f6)=b4)/9K258R+L+edSUY1[Qf9]1C
=#H0D):Ma-R(eN4^>N<AZVGP/d5;9U?-I-.fA3EXM_<@T#YJ:)-aa>VVYKK6A+.]
N]bJg(:J9VX&HTgDYKZ<=5K6#-e@A9FV=g#//Kg3)3>765:S<6eSdB(EW(@Z9b(0
ZeMKV7)9PMR.AXaWPea-);Q<(c6-Q]aC1Ya5-L5:8#7-.P5J/&LP:JZ+f)3B(0/F
a^5X0Xe[M\:1FVEK=;\1BfUb3^A@5W@7J3O+D4Bd8+=QRVMQaI7U4ZM.e(N48>b^
;G(P=5TN)^J\HD]^=OKO[TJ),<E]./O:eO9/#1W?4VKO3>C]FFM.4,.1J20<8O_C
+<I9R5-6E0_[Z+3GGN+[\@Z7G/)HS7GMX1/1Y>cX\4\1fIA[>e[[:.ZC4T\[GA?R
>_Naa#\,5T/&dc-.4B[:BgU(=@;I1#YE@fL\UU,PA7@\D5+2e<0XAd.?U@;2M:7K
AY4DF,]=MSL;BP@PLb4A)&10BdE5AZ=[cf?RIL9f4E-A5&,b4WZTc]5_KgcTQ7V?
)D9&AaY/0:SF_A]R<E1YS6>[(aW_+NXRcO.F[MAK>0ZF=G:N<-/\:J?=4,TC\WaA
E[W-FGF88)CgS5X5MR>Y:QQQd8+,)->V/<Q4+A4H2IKHgYKe<=76GS[7\\+1<_TW
(=F8.5S695VNI8YM^G)G]_XAUB6=cJIM\KMV1,OH[:D)CX=/1Wd:)g@I0JKdXO@_
G9H3[.]Z5_4Y@L;,QW]bF4&5=b?/>+CVG5S5#BO]@SG_MeG8XU\E9(e]YQPSf+?2
I?Q&&_a.=2#Z\HK6a7@O&;>HF4>#XTXSQJXcVQc9^R1RIT=]?@c9-W-MaW?1C>b;
)^=GQ#D?SCU<-d;SbFRI:dG)--bYbg27@B][f:=aF=ge_+Hb]ZKAP8D5ET(I.PB0
837TOH)^F,(K<?+GfgD/2UYacYQ5>/MI-;.@@MM\4W?(f)c/eSf>0gZ-Vc#ee1RA
>a[g=-#R.R4RC2cZ?I-&b+F448=R,)ICL78f@L\g-f/HPagb[NE]J8]QEMbe):7;
[XeK5\)bJSWZaWP9857U/P81V^N+FO_#PT6?6C(W..V1:UcU8egIW;>NCQL:&/HN
F:e_3,JRCb/KcA@@TZ0Z##EH]]g2,=UfB2^Y\>5gI]HAA))K[,4E5b4@G.PGfPQL
/L\fA=EEA1E<361RQ7RKSc<4=N,]c4_Y;gE+-6X:V0FFP^XZG1\#@Id1PBcG<T1d
=L3O?SZY>ZgBU_F+ScM)[:==09#\COENFa6HH-CJF[^9gAdXI>H)AF=Vd6HWVGKY
D6,F-2#aKZ)9Y,(T3VB]fQ3-<EP2H)W]F?d</HR9JG@cWb;S:D72N@)>7YPA_NNf
+\VW(\>&Wd:AZ43(\Jbd3fA7aA4^SS_>[3QS/?-+9e_^:9]&;N^I5TBD1WEVW;#c
=G#VW]5]?SU&.=&P7#+_DJJCO)2DKSD&.J0W#7gWX622X[P.Q/=\g:;Ve7a4\0Af
Db0^VOf4WUc-6RG]Q?\BLaQN^L12>.USHDdRNc)-g5:(NR[H14G\I@3/M,:N:ReE
QQ0::[EA;AF0_R;=S>eHOMe^Z4_dYCFX[,SG3+aLPYFS@RKS/Gg,g&PP:aB_&K]>
E9D7IOCJOR0\5e^@1L1IY-La5L#aeP_;H#Y5)4OA,Z,_#5;c(OOe4Z-C6;S6ET_c
f3Y#g9(/+b0\#NER@f&[L9LL[ZJa14ee17fM+gY1BM/CFVY]0RAQD((20C3JAW0P
#GSFM@^L\MUK12KD^(Ee-VHT8)^7JH(UFa6ZNcSHN[DC:_9>aS]2<6\Ydb6+76=[
W90H^&M+S,7BBe,IC=VL&7c-PV@))b;2M:5Z?g8FAZGM0<=cN_(.O4.Tg-E97&C4
dRLNFY][d:J)Y0f,#)b1DTI3@Ob0^/dU9&DXM,&b2,O^PCRUgJ/aKGd.V-J=@H\I
e2CWgDE:M@A7AE6(f:bb1MYRFcET<dQ7#/ZJ,7Jc/(R>8_E:>NL8:M2P\68&J>ZS
?NB]H\]K4g=VEbbOT#9&YEHdg?^[Q350b7W?.0<IRZ2\SK-RK#7@D65dAR@N?_\1
_/2/72W3=CITT(QQ=34J?DAM9IU0XDY\#6_?90,b>>;72KBY0.;NB@B/LMN@EF6>
A6fBEEbM=#7dS.HAM,T@OUI/3^4Fe_Fb?)d]\]1[g/LXNKfUCDP7a[A6cAA;3[]I
aMHFR)7]D]0bJ^>gF>b,F(DgZ8&LKX^MYA=?e(=Y1PNA3K-U+]/HE9B[3.L]YU#@
ISbW32Q#Y8Z;bdV),>(O6L;NfT?P#85K>f0b?\J-?-<:2+P>@WX#[g(0AHHZZ.+#
HZV^NgAUgTA\WXA8\b6cO,=Re][ANd6[,H-MQ4MZdO?#OSeQ[-5^LJBK<=]WRgZf
P?[eKOKP[I&X<\ObMe1,-Y2CcVAQTe..<J=D(@=.7gC5;\1f#S_O[JcF7UU.b;E=
E<\(#WAcC<LST0S,G1YL_VWWAg76b#gdRKIM^\CDg_C4&:\EQ<O]VF^(58,ZE#+F
+0R2MgaI>cdPFH)3VOJP>&ZX&^1#RBE8[MWZFTD31-(3_e&dE=08+^TP]=9HX2QJ
cD?8F<C=<ZIFg1NPS-<NN^d^eE+^RCTf/(DTJKP;fVX(?E85.P-B-Z-#cX?M.9Q0
cHc&^RI,U0=^50(W2IaCWOD^L0MQM1+T?D^UG0S^1+f0TC)@:_4[CUJ-2&Cb.(d)
GDT-b9;;SK<_E.G)W3[1F5^_V3FZ#/QVcB14I6B]YbXDYYe;;5Oe[81>P[I.;[(6
@R,FV9^#1O?_]ST^7/0?5S[JOS/)8&73HW=8UM:].>aZ@B,FXW>f5@g7C,[HK,7.
CU@.XP#_f_Bf[72UZJ;33e8/3X,=D_,&Fe9LH<I<QQ\8b@a/A/RNATP#IM]_85Bg
g+S\X-308]C7Kg>^4/LYNOHEICI;P6NKX]\HG[V8<=TUV#]AERIg0:5cE7\XgWLa
cWLK9IO2D8<3^Q)?Y2\b\&7/+Oc;UU:bg[VEA.91V5F<?FE:@:Y?T1K]:_EH;e,;
a5E:=>51E#&:eB&.KZO5+\]JIZ4_^fRc69IH0O2^IO],R@G(:CEIJfVHR:2>MJ\N
F4-09e]&4KFBJ26O<T\N2J);6Mf\AAR4,+J_NR8T=IBdXI.Z?e7ZIN16-6S#I7RF
\S\-L7;KW\&&<I,CM[a].=IAA]#=Ta4U^fL(OH.Za1&Q>SU6(&)ONdbZ9)cDKA?Q
5N/;[4_F#XSMgZ5B/dB1#g8VI5/&;XF]Bc@OWJO(1QX>Q+-Y<(IG3E;ESE<)LE#Q
,JFHf,d6#:Uc/LY_)Z,4;53QV[]]#(LdKbT\(SJQG&D\.4:?,Y&LF[&FHVMKgAGT
0g7M+4G;)Gd7]:V0,89=<C+AKWNd[#1:/>U3S)b_+\T--2F<Z;G-.ICM64d?M?ee
;G?R,#@T58J=gJ#5,=1+27+GJF2=HF@>)\6F,JaUX502<.DJ[0NB?X1<+])4;,T^
9C8R:[(48e>9=1WM>N5d937dce^3HT.&#@<(TK:<YMIdB3E.I3=,NYZM^;e&JZ8)
Q5IW@6QYeKNgdK3;_+)T>1+Sae@Q=0A4f<d=c+OBJ=2;E5D>Bb9g^Ed]X5\Ef.Cb
M\Z[A9^.,WY3?a@65HWeH<V8,/QB.<QIKY1)2g<5P8;PKM5Db\CQ+d6Q?9<]TK\N
_M(<ULea.aP&Qg,1I,^OF1,]Q/D[Y&.YNeVMReb:9N1cVJAHX-^.6_?b]QSPE<_V
(S;71SG2:IXVRQ<3B4@_f?MdU4RR(Oa9=4O949-(;3KP+OV).ga^X18ZO,>M@6,F
US9,@V\P=E3TU,C&fS:Wc8J,0YT+]JP:-,;05VY9I[Q@A0,ecPfI0F2:0;ES\S[.
B7e;IeB(Rb/Ua[@6KT1cG/9[C0&GbYR#PB95O7_L_B\.c.FMHGL95K_aV9aAX33C
&STJbP)=ZY&XBPCNNI3cTMHe;0#6FM43K@afXgg<AU6a>510W^X7J&&)YGTIKL.#
ZVfWfJ?/AX9D=RA^>B;6[L03JH+VFU;TTZcB=0@ZF\896XCbB45A4N4Z<g6JP:S@
X1LZ47XVB;9[2W)&)CKFR4(JM]GMH(OBc7>DaYJ,L[FN?B^\7\ISQ4>-<>R]K9^;
6.Ia25>c1c1-QA0aT_QYf]P4]-YGT;_65UG\T8&P:#8L1H(3ReTb^>^[8]-48Rf+
F.Bc;7M,NFB3_^8XdN;F7Wa:T5_VI.__bC=Ye&H>#F(<d7>SZedVQV?fRacW8B6Q
(3fba[b=\\_Qf.?&:T.(=bc.?..U<XZ1[6H.4/.TI0#5:S9EX5Y?5\QA75YaQ]FH
D5ZN;2(Gd:+H-@IFVad3&2\Y-EW<EWf166QXP32N9)?S<c-G_G,VPL/#)D4WSRNY
gSI2124W92#]DXVU:ZA(01>0G]B7>cGG^E?M-A69Q)[LRR)Y1S)_K+>E=&7=@bdW
,D;[b2^LFeKaaK4=C6b)SXBRAbfdb]JD&(J@UF&2T>7?(#_)dbI\;=[6(bCH=dbf
PD)d_I0^8Z&g.X.M0XgR(HJT+98-)R6G)7dKBOFNARf@&)gP(.@ba3aM5O,aOgU^
XH5&V]P)HF5d.;6+>e,TVT[S@EYI;2gM&1bB>#/.-GbJ(@9aPc;2[7PKFJN--?V<
IN\G@X\<X_VTZ=11RDUFF>E6D#T9N(QP_^@Q-W4]94;1RdSbFP+5&T?.gg6;IH\-
1:O(FbUc<JMP;IRCKE6YUEfXN70+4_W,.JLd&,FL:<XbS.Ne#aD[_653HK:^I4-g
ZECIZS,KL<)+0ZK=(@D&OS6XC+>K_I\HIc=YLA3,=d,(O4)=]03](,Q+bO(1XbGc
IEa2NH7.g_ZZM?>@Ecb/P7&&8_H#:W>GJcP^+;.fZ0/SD?Ha>][AA\3)Fa.Vd#Y<
Z^YC]f]EGZZQ@S1LbO&dDA1:.#ZBFBY>XdR)/_d--d//8<I.YGL&5f+f3Yded]X6
)S\3ZI5aBWDS7N=1F.8;cB]SPBcRNOeZ:Q(JX[0PU25O[9cQb_6+-3W5Nd:(D<5-
?f^_?H^8#@W0BTe:/EI:14EbEebb7g6O14EOf.)39<=K2/YEgVS#,Z5RWB(^Xd<\
CfJ4WB:3d/TVVEWVJ-.<:Ge>c]-S^3&O)T6+FTF3d,UDg^T_+;fPL@JB-1/SA[V/
KH?X<>[8da+:d#Bb.HHfT_R-976/5-5@]0]4OK:O)7ER=RBZTM[X2N+]gg9bW;61
O7\DS,_)A;V[1-3d_fc#A3>07MG;+FC.[+c=CS6\<L<]/\=[>(X-ADX@R)NVAcO1
Z974?C.78BY+T9J94=(E/<O0PQLeZQVIc&8BWX_MB:2:RY4DeJ<@W0&?]5BXaC#X
LN^1Hd0FTLEaK6\5=3S&-.AW4FPDB)_/MF2SF6[L;QCSMH+3N-D?&bX-+&KPg9I7
?08:ff0?N@b,GR9^UZe?GWE3[H.5gNe+5/J18FFN_F5H]cB45M@/=F=+QbLXb4(G
MO)R#b(F=&-?642UGNRXeNQ2IKPUL4KJ9>d71+MIG:cfPL,Lc?P4(T<X+,.C(MM1
-g@HFF<?0@C@K5)fSBEHMMEXVHf;=S+D16L.g+ZKZa;AXD]L,S:#,=NODE^@;FFT
(3O<3BaOW/9Y_VH(bY[RGRcX_cMS+_(:-.1V)31[3FU>_/664b9FQ_](70@<)dM/
OE@GQ@6&G&T5U\\8U3aR4S;6:/FNMcd,0[W7NR6T?A-&:2MZQ4GLK0\7Q?3@fQZZ
5K[N;3;LIAC)a&Y>)Z<fZd4C#COGbF.2P<.4N2[^aEQ.>I;cK2&UL?OWf\dge..B
?+#eYI+;&H-L77>/OdL7TBW/WMXU&IY?NITJSe[Ub6,R8@^;0>H(_:_+DfSX7KB&
7Zd<C;3EXEHB)SM5<fT\_BCgQJHUC6.-)b1-H;9K?JBIb\L-0cP@IfLUM4_>978X
cd(]AI[B#3:?=)WD?dO\<SKPK)@/O=a_?g)G(D=J-^DBO6JdSCcfR?d]S?7-&1F9
cQ?UfbJY>I#RJBH_O?=>E\;B:J/)B(==[RV;c.SZ/#NE?JOR(U1Kf7eZ](1Y_&#_
7A1;)?EU(5dG]Ef7-:2)J2(6,eY-KWOT[dcYW#eM.5a;@#^PdW8-67Mb+V6?dg.:
D2J3YB4&RfdZN3([6E9f&5]F-P-(J,#J40V4,,J/FJ4_KAWYMX:>=Ce&a77,H9N/
K2G0WaW/;]3#9S1SK47>.Yd[E].A@d95JK#93Y>)_[b=X-cGMNLee?0IJe1;0VR]
_(affSL4L=TWB)SXG)ggA\Qf>3eeELR4,L0CH-<>,a4H,O.M1T78gADH3V#\+_9)
P:5=&-I;DQ\a]Sa?27AIId4??H+E4U9C7IA[O9O=G]LF86)C;?.U+7OBHNcYBT<6
J6Z0<9[W=N11:G3bIaM/;1cXA;DJ-3)[W@EVR(T8C56?AMDf;/1O4bG4Wcf=_L19
2H1gdC[Ed1F6D#N>Cd<Ia0BFO[Q?#TBV=gVRLKRf0^2M-7SLP69+=SO_+B9PfBTg
2f3_0SdO3?:b]>W)eU;&+20HKPGL]EGTKTWJX4:Gf4W#]_3</4C(2_G:Ob,2?KN@
1Y&IQCTT>g:\9OFgHL+237J?#3T#]DF#HAOYT;(Wf+NGQBL3S[K6>RD.7UbN/N\/
<-CQ9DN0>T,6F0?#-7R(#1;8&g279T)0=H4/XL>E;6fBL(D&,77c=EaWD_#?^e3=
0OMfeU_&Wf99E?B.7MM,^^3(==<C]QIXBXcG>;^H>?cM#dUd7+RDeP^O)cBBY;:)
Mf(,QME9&?/PW6;]I9bMHH]+,?J6g.-cGW5QYS3K3P8W5P0f/P6J>bF71];K4D\d
N[IQZ+2#+C>Qb<#E.C06]1O<e,>)eZ\<70^;g#M;JWHLQ.43\K-B71d=W7H(&M4O
6M^03S/,J?EU<,Df/E400](ETYXNCS,GD-GV?Z+-\R4feY_3,,BWH6:5D:c)B6OG
<UT5M,^P]BdO_9e5Je:H.VJFYf_-gSgL<5Wec>E+C-F<9Y<#AA;&@:eg8E^]&V2Y
2Z>(P,UG2?)CJf6@4JP8[Cb;D]f2,3dCA&_K0S#G5]O>XZ=OH3?JHU]JUc(JGM=3
8<V-.[38,bK74XF]bIY[d0=9#Ofe6YU/-W,aE:7)=F5QGD2=eD)#CV2UUE5-=I8S
DQ7XGcP3<?)Kf7\C-c7^L>7QP=TJA]+HV>B/dX+P)HM;TG;#_N=5ET<@,8A=+Jd0
bZC-+EYYUbOG9((L^Y0\>-QSL@=XKI8@f;QQ<OWG\DZ</7L\6?EICJ&?T+L553>F
Y]EZV_;AQ+S-,6BPSaL/ZbbgPKA9IPBC&eD#JJ6cT?]Ye[@AXP/+EeSY]AL)QGSS
FC@MV<\F,)#=HY;J5dOWT;FN/L:FR1g^&b6gY/&/I1,+2&\YB/JW5#\U.9N7^.8d
WMLe(IL7Ad2(ZW(8(Ug)1DeA0P,-QIJVMg6(#(/e&\6QL5Xc^OC7K6_/WEXQ1F),
.(aYA8.MKAG7BE/O.^5<5eT01V.+bG(B(CDZQ(+.^@PF)Q@(FXH4EO.1J\@]KSS4
S+^7PSeFPJL#ZfGC\:6;)JDC0EA^\GJTb@05AR1WKFR4Ib<FW3CD3.;fOR6D&4\;
7>PPI0YgKLJ[_7,##R2_Q&)&.9L(H16CS4#Kf^VNH<+3U9Q[#DTQ=F13G.XFL:;E
G,&\XB3eAZ+,PY0KL1RE)_EGd./,EZ(Q6RF,B)/_OK^((^R9UQ(X?@QgWMV^[FB5
a^Ld.)[WRPc1;6VS/TOJ+aI5]fV(06Z_QE:U4:UP=MHQ-X.f\0H.[Z^C:NL/M.dE
@b8ANeJ=WZ:1.4.Zf[+OR2NMa-_[_RMH,S^S5&7_W#Q(MGeX>d\1Ie;7_U\,YHB.
(#5U#RH_7BNQ&=cKYI>e7+a=4F9=E\#4,gb\G8WFVKM2KfF&\/3;f-Za2M1G?#CK
X1gfV:11/4FZ][If^L.MBF7-J2S&-3W0?+6?.?1>fAA4D_c.FcKWA?&^NY/-I+6_
341AXOf@H,@<2Z72IE\dH6<?(E]C\9D#\J+13)(Y9G8V[2V4U0[>?<NgD;R@33QJ
eUGL_WASS28CS_W;Y&R-11Nd[\1^03&XME01+X(CbRFDMO/T)AY\0T>0#B^,I+Ua
gO;9/5)WPd?Y>I)]-95TK2O7W7dDL21RgYOX(5VaD-b6Ae)e)X^?7-35e<&:\RIL
8g86_I=1\BI\:COVdMV\RR[R>\g;8-;&9D21AQfT^@W0]A/KJEb44HISbG--G0?A
8#6E;dW=<61daL<5R9U5&f)f&VBZ(TO2Z>#+6fGRJ#^J^)a\3AHd3CbN(_1R@<.9
OU)@.;3g<@\>0R+a#9[DCL-W8Gd6)N.PbH3RbgJPE3DZC2(80#]#e:X4LJ<7T.[[
)X,8cSXG8.UZAHL.1:>;aHBaa,(0G0/e8Y.EATEF]JU4f<:VIM0XXa^/ZPGX+L38
HP(7<V/JKb+aF2_:;K,WN)[FZ8-d&<b4@#3=UK5<1X>E88QH-Tb]+5e-]]R<d3H_
S@GAD>5AXQDW[\6XGb3<]U1aD/:.DPT+D-6KfL/aa5I/F.YXE#AOR28;7#7,0d/Q
H#N<,X(V<63IV8/S34)8?T\YN6dDJ)6-JJ6f7Q#F2b,?4b\B/ec5<Kc/)E6)T66U
0W2c7G+G[,=>_7G3ZJeQ+KgEcZ2V<YJT<W]S]1/D)DUU8fHEZ49&^6[(aB;M@KGc
:If:.QOMdA?J0-[H;[Y74[1Q/O5W>)0H2P3^FB=2gFM99Z1<XaL2<)b+2N>>PW.@
f3,]fB--A[/TZcB\bbIcU5)J/\AfYIPIXQ:4f(QZ8GX<b/_8\7fU[TGedc@f-L<g
fW?J<&I(SDObR>-e,(YUS#639,g08H^Q6+2.e[&6Ud3&^D@>\8gc);Tcd])TFG+=
3OK@Ed)7+1S.4T[afLV[[7=9]1/K&]S,8JaTOgI^#;e4[5QL8^AU+2?WYP7?:K<d
8R3CQYe#RSY6:G??WWe/Q:RID-LCaDcXK+1(-UM;1OQ\7/S1&8eg1P;9a3PH;IYZ
)OL78gR]Q3^E-#MUeT2g0R^Ce@Y;3S4P(40G[\b\3#F\YH7G+#F7,FRM.[R(.5/.
G.b(b^VHX-CX],7RAgPddd7ZWe+H7+3^HUIaEdS4dA\/W6MM1J-Ob254SL=Xa,bF
&^_dQ5S[+=6L<bg8GW=).]2JE:BfHb8V\2XMC>V5S-7N^Y8)VSXF-DP@KH#I(0dJ
-,d\,;YIJb::<G7:7(#Z;U@[L;^3c[EU\8Ag65Rg<YP++J@8@Q,^@Ka_A3AZ9=6S
dTc6.CN\IP;a[(.V><N[;f_JRGfWWX;9,Q(/EXcB@1.2R/IM.RS((e95&8RV?I7,
<f2P;Ag^,XT<;MFf.2D<OJb.4_^AeIHa&ISS17-:]GCKS)OVM3@2LZ?958<B1egC
IYDRNX^TOaG-<=8(e-:c<D)WV]<<X;9#YH-#ZLPN1YN#aU2XbH0fVK2>,Lbd7Y4_
>MK<OF_[R,BG2]O\Id@ccXB86CSWB805P.F.&GZe,X=dSf-D-DQ.b@C<FCR;8)g:
NKHc\WX1f;\H51LDT8aNf)70H^?54,+cbQcAU^Gd:ZZ(<N/4&ATEe0f&>/UF5K/P
XK;1+Gc&7;<@]A?ZG^1F@E[&+f(D5)Q](JK737:#AYMM8d,K;M4fB@NLC]>5+)TT
cDO:=QAf>6V70WO>8NN1M?I6)<d2O;SQ]c<H4-,;ZSX[e4f(ga&U;]CcNJKdO<-X
ECG+;7KNU#.3/dK>@B8LU7\[)CcP(N=30fXW)H.ZDB/#PL0IQBCJQ+XP2;-M0_?8
PIPDc4D;P=caV3c3B3&U[Pdgf:2[_AV0U0^\O/ag:-\7LCIcCR7g41]WXG8;,+_?
e&F>L^R^\K5LgOCIVO/:BDgD+K@KF?D^X<EaQ+ICTb12KA4?[#+U^6d\\(GT#Jgf
P8a_)1>M]aE03Y&6\)T#eK=O0@MF7M?d8TH/(_,V&)KbH#?.PQX#U2JYY<]b56HF
K;C/2QQ<af/LX:C=gMXDV[44>ASc4/I.UfU]a^aKf\F/^/dVQQU7.@a=CE^&Ue:9
.g6&Tb@W#1UUFD\,W=^8cE@H=CF,&_G\1Z_AC,2.96<UM8#B,c&C5eRb7-TQKdLI
6IKKRNZ&c]>]]FHd\()/,E3CKXFQ516b34XO=V)e;T.B:?FSQGJY,87M(V1+3Q77
2R#Pf^I/C3NL:ARK/3fC]I?M+QO<EFcW7&XfVR-X:I[+]egegK4O?].gY3+Df7U-
J^bfOR[cg?+Y)\a4)PRZ3L+0X@(N(f-_LSII4,S_^B@?(/g#H<QQ@>#VI+>\A:V4
]W,+e/1b^7K7C[:^B[M#CRZ[2Taf5X,;IL:)YV9ZOEUZJUee@?0Cc(H^S;PJ7H_&
2cBV_>b-gB&6cLd2/-VV0.BGTY\S@22FZAVfgCgAb\94X@),.,E<ZBJN^a>)FIeE
6Nd.L+0DUH<T)gK?^d?,)A4SHT+=/-94O?U-<DaEK+#1G/NJA?7F+2>/B.X[LM&#
T<:_4^VS5e5\<7cXdY)Pd9V1<S=]Z5Y3=d\3SINbb#)f+JQK[3613MHbXVdcS1I;
VXM)YR;0)FBbIT7>P,@0cI@;6U0#@TZD#EKacH76,LM[4^H2+2:3\<3UDbeG(I-J
0\Y/WRg(>f>Y^X@MA^LX\#5)O>#AK6gM6FAI=[95K3C-,@(_ZUa<&S2BQ]3be88W
&RK5JM3(M.3879Lf1--CeYC]FTRe(MT7H9fO=g(;&,+DN&Lb0IC/Fd:,JM:W^0b1
^fM1[FE#UL:@S1(?P[)I5HB5=+V=WKGf4X4fWO?V(cC]FZHW1^?C]0#:/.5gdTER
,X^D?b^SLIc<G0#M\TZSP^A?Z5SX;Q8S)3FHJLB&#UWRK.,0)I@YLLV\MU.LFMQ,
FIe/_@Ec)TbE:HM(g:DTD/cNA+P4H]=3HcPC</<=7;Y6Jd?W(0S@7aU&eUg7_03I
B2EV8UO30?TB+4eWPHLT[[V61]R.=0\NedH-]a^K&SM5+fb@-_1W3B&DCM7_]>)@
bR^fWZ;[Q=,P,f,^SA57Q09U>&(;#KX9,PFK,#bgO/WPd>+6Q-/E<V(,7-&e>U:E
JV716;E^G-Ld#SZ>P&.f6aLCO,Z@GJK9LKV5]OC>)=-Y6c4(@=&7CA7L>MWSZX:6
=U;J-:M4D25V8:fHES-;(9\7Zb=NUaC.@]\=+^>4,&NFVW@24/A+G@^NZ0<(TE#c
EDZ)UTV[W7?M/QEZ,];Ga:1VZ<XO<CE2NPgfAU9S.RHT&M9@L0HXfEW9EcK:[Qa>
)#>._\U<L]F/Mg7T.3^Z&f\F6^#395T:,0&[[<.1M81^cWLJV<U8-S00[\5]:.D2
1_#HT//^Z#D0(5R,XK[^Z_\-&D6&VM-58E&MAYG3P-B>M/T0bM@E:Y/W^<3L>4#^
=UWM;U(P9O<^/)_e[gfDNI?.Q]b\8Y[f<c?K8YROe8MZ7a6,a<;<,A.Y-/WUV&fK
aGCd^?7:PQMOL9,:2WG8PZ:2<]OQbD,Q)VfUKU\5&F37QQ/FM1[VCK9^F#efL-U=
fF>X1V3FbN(g2cC1H/UBM#0I>&NBGe7]f\/L@Icf6MPY60(F5ZW@16LS,0]@0fae
5:?\^60.3D.b<e))OaG#Q^/L.-HEV-DCW>L]Ia69XNP3S.EOGc8eP491W6-]Qc:5
NZ+1FWaGVH=7\E56#BZ4>VFJTMX>01_N7X6])VTTRPcEGGaE6S1-1XM;)X@S,IZ4
>-e,PL=gL[cYg[D7?^LM7Z5V^LNKJ,fcUM,Be]aF3C_54F[CL5_C20]EfNKH_NNL
8OA#K)/Q^.CRRe[-Z.[XF]4Sd_VJES]Z0IP.fb,>[UX\KgY:+@3GdXDM<=7\4bLb
1KO]X&JQZ7?M26_TcRMG1Y>e<T=;6@CV)(NVM]X@XEL(<:/ORA-c[=[([D@F9D+N
0]2]0Z.VB/K?LP.EI;^Y3]2M3ffDfA+2D_=E&W][A)dCKN]Sb(_#GX2gW\DgCGKB
cFOQ9(;_d4ZN,6bOe=FV^d;2#dfF..U0/#W#XcM?Q/fbJFD\TIZA4?=()(+=M/7;
0;f8(7[JY,8(F&.0H1\FYK_Ne3MRAaSB9HgL2ED?J^=a>-][>>B\DN46.N6:[T2>
(HWR2F7BT^M((8f\d6Vf\ICG1.4.5S;N/PZc-c?))6J[.5J_16QMG_0Fe]5,gTR9
60G:cTJa)Z\CNX1-PIc_Z;5Z1,G7K.._U[K,G:J(b#9OAKc#74FN=H^X)>2[XTDT
)&-&_KOZeVL7bOWUg9V/-CZb(K>8#PUF^X)?Z(8,DC,+O6DOSDeBKQQf>-#88a4J
)>59-QEYc&bOH7\8RG]>ZF(;fW2a<D>:g[UUQEERQ7V^MB^F1,LZ;-V(D4#RNcP_
FSc0c.ScENLY/B=;\GW)B+K@YVGYO.-HQ[:A8Q8^^&,-O0aKUF5EVLO^E2YC6++^
D;;WH8,@,O7Y1R8C)YFFLC##TAbb][\U6IITP#EcSX[OGTD0c&FW/=WaF0VY@55]
X40HOaQ/O=0VPKF3A<>=QVbETY9f?PC8TQ,b12@aQSDKgAJR0CEG_fY,XUA>3^FY
E.\g>;JDQI-Ma0U#^+7;PV^:3Lf&GHYRXHAC?=7#WOA]6A7[=46L[\R(&QaRY[5R
U.YBdJ?)IQJcGFHQMG7/7Y:P,,Gc2c,B=7>K<RMA;ON81:WfaCOHe)eVFR#8HN&X
-/=6?+GO.?^Y>ed<aFZ5&954a)F/;4V-FF]4T\[4f8RW6U[AO8(?a:d@+4;[=-K-
gH\)]&g_)[)C8;W#B>Q+9Ng/F+\U>K0;RP8GD5bM)XB>C4=Me=R&WEOGLY?=3>,:
d#&U(&bDU+0E[M^cM=IHV#SB<&6e,)g6R]EE9BM@7-M0&\M?8:.@X?5FNSO2b.TO
XCX8d5KOBC9^C6bSQd<5LB?3Hg1-N#(L[1#K=KU4<)4H5F3_-eW>/F.:KT,LEW[F
cE5,MIML-1VcUb(d8P7FT=+W#&AgG,23f#T&=OJ2JNb_F)Hg/T@1L[3#S(QJ2Kc@
4;_PNFR;W@GHbFCJ5#4?6V1S7>AC6EZN_F>SIF.:@KV06g>FLX6VSe:MccY+2_&g
MUcJ]H&V^Be;^=EFZT03H7]_d>\-JFV^V>6J5TNE>#d,@3A1Z:HH7A@fD&U.WXZW
<ZLP^[^c._7?d>N?H4WO]L=]1VMR35NQ@6\;f@^3>-55F\5GMU/Q/fMZ4U0\-QCQ
815Uf5.&&G??dXR7aVASFJSA+gf[KK4/QaLL+7HG+:EaQV,R716ac6-_S^>?VMdR
LTH->VEZPZ3d7J.BL<<05.6W]&/@SVTGX@ZDV5B)37)=5;8>B:/g4Z1GKJZHggXP
LU@@)6L?63_9=I-TTUVR3L=E&9HEC;W4Z0DVAHFY4J/UG8CRdBU/+4H5)JTESE#1
=3d>O_[+I]ab/?^;@]V@U-:OeR<f+6g)IG0>5RM2/DOJ;IVCH/T;+e[gLPe;O]aY
V5>-]M7fIUW<:MB;)S81/<>O\-,NV>7B4K5Tb=_76U^b6BYH]Ld_6?2O\-.);-,7
MM_D7)a_Tb72bRB8g9##UAE&f?NW8a<cQPR@+P:fT:@G#SLVeb;KDK)dgbJ(J=X=
O_[_;9?D1Ub@WHL8fSg+5M#OTSbO8AfZE#S-)>;UTU8I2YX(=fBT+:1#XM,=1&>S
KCNe/fC&:NYC0EN\/Y6D4gQ686A+>_Pb&O6(W9;(X[P1U0[S9&?ZFNUKcL]@953f
.J7ST)M1FN/:=0c#>[M<=U0P#ACKKPe=J7&@ae)[/NEF)\:d^)LJY=N>G>+fI&M[
M)b[B0Me^>/,/_;;EcUEKLTFPA_ND3O#K.5QgRS36cEMf0@^:A#a;F/bCY2&RX^9
bLEb&a/)6,b.-UO-[/QI?+A_c(G,S7)SXW(?.^E,DO7@ZcfYNNSX5+(OGFG<-/Ja
8Z[V/VHKSLJ-OZ?[@6:MgV6;G=.H+,_<9CHAZ1X^Q&e<AdHRS.X\V0A6[[@?Q2R[
2g-.eU/Q9:c/-7V,WRSP+G\15K=\bCLXXV7K)5DBK5Me1cD3d1A<OH2S=/S3<(cf
3Q0a[H-@ZYPPa&Q[AG:g#^(N4G;9E5fc8\[19,.>.Q;/Q4RVL2GTW&E;QJ)^L#(+
(?d4E41NS61@RW9Z,GF?CL8TU-Ve-+F]].f:O2Kd<<HDe7aP2N_J<#]XZF-G#T=<
K:b@\\INLIfAE4GW=].82#YS0ZS(Bf0<0O[?PVGZE@]H-]KQ<gEOWaR<\]+=&FEG
fbf?ZdfIZ-UJ+(SB=)B9e]G][==;Y/eL>2Y:d&UE_1\N?M0g6>58,FCVH+=&OYW#
RDSA@WY<#T^W8=N/Q9R81E<4O5aP28=\NJY6=fP;N\9LSN10a7-8Q)A)XYJ_/X\N
g4X,LG3]Xd1Z,92.+[E^Qb\R=dc2&+.G8UU<=H6Af\R=L,_<cg4IQNQ=\C>Vd6F[
7EN;d<g4-O4@BRDE#4PX171H]NC\_U_P+d&<0X@aeXQ@XRN>(=\]T<?3BR#1Ab8)
#BZCUC/#aeF2T73QQ2[a_\^(+)edY5=EK[HcbPCfZ+>b\e<=0K2VX1cVSgE]TLX^
]3)1LYU]]aP7S4I98B&fFDG[Gf_J,X\XN.=:c1e@_05[M[BI3S+^bfEB.9KZcE.9
J0^2SLBUP7ZTWUb_=T>d@T7T9<[C+J;JYgL_V377R8DVD8)3;GMZ=N(W_+Q^/UG2
@WfMB6SEZ5@U#STZRV0[=;f;E@D7P_FRdFB-@3/R_/]c,?f&XQ5Gd/?P>J5R)C)g
MHd;2d4e)Nd>X@e/XLHJEg-;dFP9cY1D7D[M5Q,)O(NA>fZ&Wg.G3c1[6>(8425/
T;R5a)?9VMWGS)2NMT[.>SG?)F\+UP.1V4)..HR_AY;9V]=KD#H8BQHcWa9>818N
DOgU2,50MJ#B)(D-BD/\S4]bFGa9cR&KHC2627dE#01B&14N2OM]HX2@d1a-->]Q
V(g1QVTN=da&P:RB.F1;;?&QNR3&PF@Z^OLO?S?SQH98S2ZSYF#4N.1a2f2d;)>g
N0g1@aP3[5S1CEQVO-@9&BWR,SWXALRN2?-QN)dKGVQIK:b6;+P0-f7;16XTd(]_
PIb/IaQJ[S25?GRfBPK<))4ZBG9eF67TV?<ZF:W#,;S-0Y4;Le+U9c45.VTLSU/8
TYF>Z\E+U1+XU=6]..\RWa9YC#7gdQIfL-3,a>3D6R?:^<8U^Y2Qe;&BQEDB>UfT
2SA9K4@I)fG7Z@KdE_P(,\aPD5ONJFG+.VNg+F/Me-W<[^)-^YCA9H\7d;7E9[@c
ST1VZIU6R\ZKI4EQMIc_<VXLgGP>5@M^>^U\,70A9T)g<R,Z.]C>(X__QP\U[\=;
5?GO<DF.J5Mc,(CUP.XRf]fN]<QOU&0\MRT0Z_D3IS<73OYTQaDH#dNVeMVQ,T?g
#0a6RdeW-QMNY+E1Z2/=6FBaDI1(>32MFN\Xb3JA6#7HPJ6O4E=QQ<RbTDRaEU[Y
L-Ubbb+5MbGY;FgV:<T_@L@I5CB9?e]708SV\A0/]K6FF\Mbb37AMHO>YLWR^8>W
=c-E5/;c1GEYB\a7U&V(Z+HRKJM[5.M>Q+7&4;:N\ZT4PJdH3Ya5g;W[#^^O&H/a
bP628]60;]S:QURWM0Z3Q]]A5Nf&S)A?IV95=^M1]+5BREGVX8KSO<Q2Y630U4_?
O3X:CL;@F;B;@E8D0GBWHL1N3[SRNG6(cAGHQUG(BHg[8O]W.U=,cXR[[/HgJ0,f
L2E^#X]9DKYe\I,B8964Z^TLB]1-5WYP8=)JMGR04Na,]1gF\fPW>g\N3K\9PY7_
F1&P.\1VU-BR)9aaa]6F29^]>ZY2:@ZdOeda88/Y=/RHQ?Lf#^L2cV(G:(WQ82@E
LYA86OSVcHUNaAbUL=^d/dCEbPUcR<>@XP0YXCSJV\FSO@RD-1g=KS4JU3;Cc@Z_
CPF8G)TBB.:)80^:TI6&8@fZ,NYP^bN,)9-.G5U8.I>eW?RFXRaWS<,ZJUZ+6YZ9
>/3T5J?..a\.Z4a+,?,?3]X3A1<Hd14\>+D6,0g<KR?QfN/VM0f1)\25&57?d1:H
^D36N]/67.2P4(O2#R:g;=>ZSF-EAU(UN0>7]d6XE79.BXB>cbT7T;&8_Y6D?MOB
[ScNaVOf,[bdBc8U0J0B0J4SD2#EUa)S.;8;@Y0f&K7c>(A5[_W]N6bg+,NLWb8E
T[b2)47&6R^@I?8XS57d3[1Q/34IP0O@cR(G(?bc>P87e-cWO0+20K][&,PaTP&7
_/+@bF:)(f_D?N,H0QC+R979)WWMMF99BGYGd-#?9456?b]W&d=C\SS-F9LC<V/G
2^581\#;>Rd_PZ>-=FM<BCZg8Z<_MP-aA+cceIf\eQPd9B/a3L(E;[OTcRN><=C4
e5/&/K]5X([+6bC]K6PDd/C67B?f[BWDMbf0=,_<IbLQ)X8Id:U3SP<_]T,:fYMJ
a,.15<f@/D5<J_(R&D8+7<8.:(:0g83G)VQ#J7#OAQ:WOKAUX--(:V1Kf(7F]>[U
K>a\+a4-Zg,(-XXa.LfY].5Q4IV^2Bg&&gXXEcJ<4:1UVC1.GFMME.<B4:[^-?NN
NegG:3@]WAF^[gPe.:b-Q9:@+]/AI+ISI-a;b]\7+PB4FJP=[T#A8PX8W]efGP:2
7aGB[UL5\fe&g5H[(Q5f9TA-7JGF3JH.Q7D=^X8UL]#\,SbV=DL,H2&0D_A]7>YO
.33U?J=6DRG/QNBDTf2?cB#)+/J8@)CI?M6.SX<Rg<]&R;Yf1A+,>UQ^9c/LB.G@
HWQ.eX)06]4E<)BCU0<^SUTAODANZKaV2\OL+Mg:)Ie,>FR4MR?NP;[2,..N(,L1
C2<Q=GDE(KcaF6b7QL\e3#F.)-/ZZe+.6^L&XY84RfgDV0C]ZXF[B=3d>DY2b=XY
E5JVQ(f/faNddPXGM@4a9Z^,]-L),1NC24HVfOI/>8J6K[bP9S<^I(TL@A=K=:UX
^M2;U(>L^(f1WPP7O\<?7E+_PB4\4Q:N/9?)UMGIAcB72bDV9\)JP6.d+8;LaG<L
<@TaQBP7=&P_RJ=WYRX\FMH7?9[5\6RTFBO/b?97\>eCgH,d:)1>DWaW<AJE3M5g
N0Q.ae:9Q07=PZD1F69=\e2d]<TV13H/_ZG_7L>bUa>b.G-;?DYO_H^)?>ZP+)1N
Sg5<01-cH7WFK4;(/TU,<T-b<)EBQagT;a_B8YbW&LKfV#X&/OHBU]1XZ8GgZ8OE
6(b,)3J+_#M]8B+Y3?Ha[WM#+Bf3D::3&<CGbaEQ#@.E6-;E3Y\+fQd,ed0QcQ^G
LfV]K2ZPd2RG@Zgd?7@:\9P>7NO=)f/Fd7Hf#]6\^DJ.46VL#D=G5=aS9@3G;6B-
XDJT#4N4e?\H<AIRO2F0,e<)V[7;<XBT;]NWTU;AEfA==4M-g+dZ:_+&5WFLV.S7
F5@_Y\ZNc3bZIFW,PRG9&dRXEaUJD9.#Te288(>W>40GEC3_faECM-dIfB?ELS[V
3V^8=;Y9Z82e:)(Q_1C67S+d:R9>RXaB3:W<O:EU^)?KF7IGKa18&M8O@4.W\7_P
+eYcf-Z4)cZ8c,UA48Ia)]YELb(Pb;_Z3LG6b5&Y1/Q;eJ=2XEZ/.b<U76BP]^35
=O\9_B^Z3[(-BP]M3^WLI94Z;UaePZ+c_T:LE#;<9,e(2YS:6XF_ZFSZ(WaVCZH(
+B#L;YL23QB]GS5\e7#QOW^a8e3[0#a8b;9TT9+&RU<Q/PX8e1>)Sd>fT44Qc6CE
F[3UOCW7bCT:X+4G]ceG3Q2?_C?##MSE^c&W>&7JeF-7]5]<[)SOB5R/,9Q2G8;3
G,g=H?)+cSPFT.T/(>ac^9.A2:[8LCJ<&T?O&\74@JK#3<Rf[5V_K,ZHc05O85.7
\FeO609=^5,^TL;XQEQL#3EW^80;QOG4CG]RWWN\\3TKC?N.R^-JeSa+Y[XG@=X3
Q<(#7(Ce]ebcd@<GCT#8DOT2;RC0V<JB1.)\,D2a[DJ5L(8HMXFG<T:.Z-aV>I1+
&E>g9]2JObHgF<(@V/R/.4FeMfGZ+ECT9>LKd7a]JH;#I8/^F5?:>GgAV96PO6E[
JPNR]BTfWQg)cVgdS9[Gd]b^B.(#S/1:6F:+65WC-5I.87HZPI;O-YMcCZ?F5<&)
a\58SEgb5.ASI_KKO30D6\Of7#65C&LSc9#Kb?8X7d3cH=SO5:6WJX9a=F3f\HVd
E\89fVK<c[@e+6R6EKOV(\XM?7eAeZ9?45[TGV29CWHGS1C8&>;?#g]W]Fd?LgMI
(aD^1ZAG.[?B4JQ=M)AP0:FY9)4V:LQH&O#EeE7-DfV6\@D(W>#D\M.50G/-g_e-
);[cR4Z5/J;Xd,b<g66F,GHX.0.5_SF:I=X7WKAb;=M2SV]gWT4=cPB7G8WKP\?c
47SJD^JaBDU7/2(_4:L4FDd2<;0WKbG?CZV7#)X@+O&6TJf8dY&S?LUZJ,OA&9PC
AgFd#:WT/]8.HSUQE7,ILG_I>#H3?Pe596Cb[gBVKaZe4UK)Y;M2cIA4AC##J0bJ
+CDLIMgb4\B.8&_U347_Qg7eDYDIZ\BW):W\Uce&X6A#TFAV)+]Q5M?TECRB[=_S
=1V6-P;<]fS.adWR@MaVPe9Z/>UZM5=-F_HI..E3TS[?T\0SdT=:/UDdV/NO2//M
3B>J/W_=..b824PLE)2FU=TfE4aUb&SgJ?_0RTPECM]P_^W2Y&dYZVXdKR+F3cST
D-KL<G(#K-EWY(_<I(g+dQ-W+^><=J41OOd0QIcUPG1VKd\@>+=7<gU1F#PEUb2@
5ED45T>-MN8c>Q0DIA#I.-T3,/4=bGM+\W0=R[MH4Xa#G(K+2/8[<BgNRW41Y\^#
#G4.>14V]U[@.cTV<>/e3O8aeO4R#ZK2X17&/WST&C,a-?Y\AH[SB>^A@3,>JdN8
ZNKB@:P#N\\OW+/6XD.)d5?W9PA+;?G?dB?(+W,E\6J6U<86@/UX7/B=<^F[GV-4
,=90Qa:edZf0C#+7&R0&e,2V:aUAWbNE@Cg7_=HXP^2,eGC)TbSaFTN@MdH^5:aG
I3+.VT1Q21-]2#F>2)(MMN96KQEXTc<IQDeGK6A:<S@gNZ+L+;&J6,gALaHR;4dX
eXgW/(5/D-;;+EH^eJ).9<7cd1-F=Af>,;9]/#b]Y(4CQGD3McIcJ=MA;a+HL)>3
NdO8EWM-aP(>_<X5e0P01\1)e]H1P44DG.UfFV2A4&9Bg81#9GcO:01^1O7;W^KJ
+/0bebV;E&IZS=V3QM=2H1#,>O=Y0RS0-2-/M##AfeAXgG0eS9RQX;LVPU?@G]9a
U]AY#QUDM@M&d9b()8QKg#N5f]X66@:@_#,,;b;Z@3^[V32\T/&Kb[[@dX.T?R8b
-c-c[-^W:9T+R_ENdcN<C38GbI;@8+8AWB#G66I=W#-#3,FeMd>T._Se?5C>dA.J
4I,>MMDA;)^OJVLV1b?8eB4M9>MVL#,5N&5LRLVg?D)?5=a5J8M\JZA<N6)4AVZ(
cM<O#_X?=F1D\NQ#a4^P?=983T,D]2KV2<T/_+9de8)<:P>7H\]\#E&,CIT])BI?
[_FV6FSB[+)#V\2Vb]-&&E=\ND>=T3deYX-a_L2)Q9KfbbWE]RL^KKB[NZ2<?_CC
30Q(1+5WSVW&T#T#,.WZeFR32K86d;:cLDA1ZPVP@>\L09:,e0UNB:Jd@.Y.+FHE
7C/]=72FB/4U^dF>9@NOH#^W3KN06ZD;eb1#<F^Rb>4FF#DV,(;;+Gg;)B2#YS/=
-62&c\_PR31#RBGAHQB7HLNBY<B[9JQKID4I[fZJWbb0b?A?Z0A.WKBYUN&[g9\/
9C6;\3WS.DAJRX(08O38E?Z\;+XTW3C)@e_F9eY.O4V5bG./YFg2@>2299;C5\>0
WgY:BE5\c,T=E(P]cZ(L(6cM2K:DH]JA5eIV]XOK&EQ/PR0)>3[W)IRJd\:U\9SR
ER#@S[Q2^.KfI=U0?K?ZK3V@KUcWC-&SQZH[[USbW[2e>R@=WS]WUX@+Q:HV<F2@
Z#e=-A69-bba2bDDK^eV)b4IWHcg6IH)Y2YQ5\]f[;a1>cMNa:.-RWH><d9&gaZ\
QIJRc6aK7f^S+gH1,O<HM\Y=A?_VN,[S2S0+4a)AdQEI?[:3JA;GYNXFKOM=5/MM
_\F<>P,F._<?=[c1Sbb81F.VGgE4e]HE8d_)OZ.(C-RI+eZ4VV<[[a&.T>JD@=81
/YY1\T.EZN_)1_?(S,JW^aPOe0(CX[^X>C_SDHFNH8[=D4<-_(dAbQW1JG:2XW)#
IV>F]F(6EN(9\(YMeP_ALW:V)D-D)Ng29BS>cJb7YMag+JI,,9.]0:&44fDV9C@:
M]AbIR05GY#L/_H_63Sd2c__#c&/>[<HB+52G;JQ9BD,:5^(gV[IZA7U0.RWRd/Z
B+BgF)H,JL:WP8LcZHRDS+XC+8/ZHV5UY5M@G?=bTb9[>f^5O_d[fHL8/4C<I(&7
.DQbcT-@HD+V=(:0\>6WaS;,H&C3+[7eQ7a#JE1].d5O#\U&PVcB1[:U?KL7)@3@
1.g#;3;CcJb>K=/e5KNCf>d94MILQL[_PFD-S&CIL6W8BB^&GS&^?:e?8E1F;2f(
5:=2_&5dMS@_1PC\Q(b&D><[O/-##]J35WOZWYE1LbUSbFVce;_BJ.X.95:Q;X_3
0V0dOOXZK(F>[=4bZbg+W81.((=R=40:8#9Df/L2<b)V<N7PI9\>U^=U^@7>1CLG
JE7T63-F?W1GLg6CW3b=bG0If83,2HXc.2O;GEK(cY<K98>_D\=S<IYFE[IGMCg#
GS0K+AH#,13HX)4?LE/5J5\P#(;WT8+D=5Y3HUdBDNcB[S5a0OX_KPVN3(,7AFgY
1a\;<dgE=Z>RaeGK83>;5P.e:bfYPgcQ>M607@@(0P1>D=U,U7K(-(68Ug\B1bQ=
7^7R5,)7[<#Jg;)32IIJU[ID70N759+<\HBVZP5K(a-L4.[fO@CQB0KOO,^c>a6P
+D0HQ;\fbd36gB.a=e\,[fDFZ\N[,P?U]I,>H^>=]N0-B<c#HJ]BS#\dW&L[<H,N
-R0gWXQDcNB&U#Wa#I4[]#7f,J((UF^[PM#f)dM8LTB;B?@<Y1)<O^6=EG.GSId?
;0S8d8L3e2-^g475Td\XO(?FeDLbEXL,AL1&&b2F5]?D?f\IV]X.V>[(dZ)]R_\J
HLF#T=7N[^E(1EF3Y@&Ma>#V\@,K41QYf:Y1X7:(&A8=R,ERWJ#@3@a1MY2;5eQO
AaL,cR=22:CZ]bZ##=Z@Pa_a:,6P3&TfNQ8(c^eCB957aJa[Db6773d[CN,RDZ0e
1SQ(=H#4Z20(eHHP-68NOdY.0C3_A&+9&.X+XC1,G6CL+:#9S:OSMecZ<2A06GaN
]cB09N:e^.]caANdb?E<_;L_27)59A9a14ET)&ODc5A725AVc3ON4]Lga^.d,]8V
Mb-dR=U2[T6)O(_d@1]M0GUgP1b1d:YgTSY#A>1Q[9M+)BGLC@FeU1Y&1LF^CWc[
/>7O&V&(^WG[[WHG8gCR1PHXM?K+M//1OW>T;4M_GA5VJ_2DPTL<U-d1BdMT[-F:
\:DI[G[AG3,9]L@(,g4UAS<W,TM@f#aC\-W,U&,]7b)fbCcBEc.J1Jcg.4#)+JeJ
<H=]C(L7eT^MTRb?YgP7/?\TaJ)&(N0Z.dMG:_8K=;fd@EYB)W(T04ZN=00\E?8U
6UWe\#YJ;6YZ^YN0&X_R^BIK+bHD==9GRc\51AQM+J@<#a4/Yb-#&+69T)07U+&&
8S3I^9>,SXXN9<A=QbdY8B/@(MF[DII-b)GaUF3>OU&HIL;6fg?0B/]P/SfY[838
5M[-bR#Tc;f=WU8OU[9e=539Bf2__fS0DRTBcX^X3T170BVdWE[H,cHZ==LWASP+
P7;V_M;7Na^4A+8J@KIccfU/NH-1RCLL]O#MYfV]7d,?9AJ<?&eb>\6TE0327eFF
I#f_QK^UK&5:5Y,R:IAQ/fA;#(#X2DVbR.//YBZTCBJ2[Yfda6SCVQ<NU1E4bF9Y
GYG5AJUbE,cO4(@C<\C4M/5e<5ITQA7EF?&0g?K_+SZ<<SA@/)K<+1Z]B5/(T400
]f2FJ)5F>IWd3N9,OBVB=#TV-D^<&bEPXdPe9bD95&NRdPEJ6cY?cJ\0ZW73#c>)
R<0=XHf[#^Jf2P6gdF4U<33I_]D<?>=HF<=PS&+ZOH=?MV/_##IPV-EG8O6:3]2/
KYKaJK4>aacXH7NN0GP+/MM=B[cdOTbZ&eM+bP72#EY.FVad-ZHbQ5;5D85WO@LG
BWdWH[,J9Z:-JQPA7AL34T?&.Ya;EF_,>Zc9=GXD4[LOL:PPN-D30([KQfGHM0:?
9QA:)[I)9D?WcXTb8-d/YY;+\)>=2BSgY8I2SaP8A9<OQG\KTLN>:&:D,;8XA0U(
>bFVP\?gMYK-;Md#1(-=#;Q0/5SAMGIX&1>Z<R@NP0c]X6dW;NSYMUVEfCL;JEW-
]F),D()1)#<]/C:UX49(?;O:GKYK+X]BQG\[SIN4/9[Q\T-YaD;0D0ZU+NNEDZ]U
M]D(PBN+)fW<PEPcQ5-2K@9])^[H)V/,)4V832Z)1GAV72^LGd:E]<=dfcVML#bc
/da-Qe,)]b)&(#)INWgR&?B>HK32PEdeRFXX.Qb,9OGfX1e4L0CN2-Ma)&fRKXJI
<HcHZGN:OZEBYT53@cN2I;Q0Dd&VcSf:OA:,ZM4?9AgYcRI>dFF5X+J+[?-M->SH
&85(LJ@T]]VgF^df;X<[PRD<X^25[fWLdE0<PQIBY?#[F2RU24@d??.XAR,e[Qc9
A\HA6:R)J[b]ZEYc&EEUQegS+g(E0#KdSGUW,0;F3VfTDRQB?ZD=@B(-4fA0.F,/
K[IKO]DZZHO1-@\M@U1G@:Z18a@bD]c/:10,#)QZVEFJ]927;38Z80O;RDHO_C;<
#0^DLPcY7Q,[/G\e,cf)\^5Ve&+(24,C3CF4AYb_U,d4eb):T.E>[<(a1IaeV>?B
_cQLT9#=ENVLP#+@)gMRT/fCIg#8E_&8^8ZMDLD4ff62WQF)G_MM]0c^V__7d<&A
57=V;Tc?ZN(dB3;ZBf<Y^OM?M=N3/T61>]\,1B.G<8(^XM13=e/FDCEDG^_IL,N+
K<KIX7980gUDP\NSa]Q.]EUL&YYZN<O83)V)e-fH>P,[KE__N9_AFOF5fT17g2\A
Y/G;-:V2?;c[eJdb?DQV+gcIW^)O-68bgE,>,9PVTL&FQgG>-9fb(B.4CNSGPB<_
(312YPIAFd&QFA>A<IKS4/:c9,XDSAZT5,_SgMX(19I?B-B?B^H.<MNA#K5=eRN+
L@<A;M_eJ]d36\:?X^=PAR5^FQ=;?<)Sga+3:M<,+V<Q.D\?F?cF8dS?;;5EEY(@
#9V-FfS>4(SObcV-,QYCD]>Q][?HP.8D5:FS;6G]g(D94GJ61PQPXL;K_;(gIE-U
W]BDH6ON&]J+1DC-BcKa,c17F2@W4GJMT]U\L?Hfb2a>/f=16(4T.gaGddR/8FLd
>-OgF-F>0M1D.XP<_fOZ[3UX?W[U&B+KMX)YP[NeCRQbUTH;T.T;)8G2HO)eHWG]
Kb-SG)FHFU)g\FUZ]QIQd^>gE>8,L&8XTE^JM>8CZT(JX)(8N-4@C/@P)P.?&<S\
(cDN#ccJU=;F3^:=E5:BJ&bX>^JP..-H09c@0YDOeA/S&8<#a2,&bHXX>Q;cBCd,
K0[P5-,Q_HKE^a>/daf;DK=YHF[R2+b6GgO;E?,RKHG7:0>MPB-7fK?:&W:E+FDV
T0_<W0C1HK:VA(C6I7M0U<5.HZf8\MZ.+M9-X5A&2,_O:/?1L#GZP\6-HY)DGKc^
7ME/g[/BB&5<fM\e?=BMY19Y[E(32TQSHIY1HV=G/59e6?a:=:G?.c<G2Z3Wd:=J
7R\A28bTT&dfL;[&P:6F\]>0Q1&<QR9(F0)AJ;&+P>Y2@5a;_1;1:H^-OR0.XgQ?
S4_2:_>&>JbgT&WReWP[.3g)S4c1YVOgVO/c/[:DgcE??[<8C_9F-D,U,IHYT/::
e=f\BM)Z&OX]=Q^?=^f@Mb.R+3(O/>&EAYBgI_F0MN5.BgS:8/6_..,C+642;b/5
fE+H4JG3>(3N\cQ_H/T3A/^C/4YF(]8#E92T_XQ=dB:\BD7BIEJ>=F3VeZYcMB8K
KKTBI_+ce+_&:/+^OROGJWT2W3EM9Bgb9ETGCBOUf?P?fD<F)7SLW4.Yd61[gVC?
IAc\(MD6FcM8Lc9V\I>3Y^TBTZ0C],JEKUHFaaK?]DA9cTY+Sa&]_DG8_L+GcR^_
cBeg5G0a-]S_+_HT.?L>?42ca<&JW:_.@2)PH-5BG;&18NTWT/LRG5--3@:L17VO
LWdBe+@#3Rb5/V@OPcbZ?P;aX[M(_;Pc^/:,=@EKe?-T#S?,0PgU7OG[?[fU/PDE
MgIW(HM+J@5T3:5f1&21.?A5]M?c@FX>cZ,(6fcPIE0e,:Q,TE[gW\0=W39J:R0]
T6d2\f>cPW:GDFYNg>66<><Q:5XBB:g=4\D\]QKV]#Y3F,De/QNIbG)@_@ZEWE,\
IJE@&O[6>9PZR-:dVZRXC-01d\7=FKT<g9fWW/]/eOG<?OPL_VODD#]XQ_b?7B&4
\e22HA-7GQfQ\QV&]Gf;UR6>>ZIHT:HFDe7P1(b&gT[_c(8E2Z[O[4P-0FfX-=1U
T,^[AM[LKYRc30,E5U;F6Ie0L)P?V7@6Jg5g:[bDUP?A#?5>aQM=U+_YEC3ROS2B
.EE6))d[,U^>AcE@JRF4gG7/P<Vc7LQA&5PB90>3a6[8\#R<^BF8PB9;:.2deZ8L
3Q1BNUOaGF\.63/Rd8[(<&=bHA_C;:&;B8/VV6b+Q[-,;f\+aBaOKJXBAW#SOI;N
\RY#ZPH^-9@<4>SO\1^O[<e>Bb1U\b;EJQQ>I(]:];RH<9_b[2(f#77D0Z<2cJ6J
H7+Q5H5>(19E?,X_Q0CKB@T3(G4029;KZQ.L/fWT\ag3:Fg.^cLAf@gK?>6[e=]J
AgOPAg[7:G<fGbW:_EXa7GE@KN(Q1?,0964ee=4d^&X,S?.cQBZ3V@]=67[<)B)L
4WJW>-Z&<I8C#WabU[bYSB8PPYg,CCU#Ld33W/]Ha-V^P-:;UeMN[T4FA=Y;1g4X
9A3JdTVLU2MRFAYgU]L,TbK&eS(/?14H[XA\]>CI>bI(]3W-8-XVC<_G#NF80YI.
VMaG[4\cWAbVDQZ+_97+P..20]W(BX<[4OCa#F.(HQ+-H0L#RE/]HO]X\&fRM@WT
1>P0O7]GS7JLbKF:U=-NgK<<1)UKV.;6(f)0]E-fbBXdg.QA\09T41-D<C5,^Q45
])6Cc0RD/=e2[dS>1XNgG8Y05?0I64]=((Aa4e/-:c[.SX0Y,eR7QRTLe&8U(>:[
#YO)2ZQ?ac,]0AIT9E:8[W4dQGc.(#:\aE:0F]H()L2I))0?fPOf-0aR:IIW.Z>?
1Tg3+UB9IZ_MS@^>efNFcBFc>@^X0;]P9OI<f)+95EfP_;@5(48/DU#G8Vbc(cZK
6UO<:?OCcbfcc)7AS]C+QX2[;N.[;?57O0(g9P>2e&P6SGALU9d>,CI(b(IAV-FI
TEVE,<+a1M,@Bd@MW/&&4H2^(dP9-FH>-5Tb>S/+NBN39^M5f5+M^_#[g5)Z6-QV
;E;(\HG-;7dQ(HQQ(H6cCXULH?BOb3BV6#JL_b,QM7U6R]P8#7O4.6)^QPIM2WdC
+J+)O1E\2/Dce4.,_1ZP5B@a?Vb>GLE5HTALfF8@WAa\Z].U\V4LV=Ae)MU?GJ;@
BMf_CQWJ@#XE+a6&Gg=a&&M:YOUec1CS0,CU&Vd/,=.M65cKH^ET=0/f>,KC4EI\
NOJGcL@QOWIf\)-^<B.g4OS,BX\OAN876N,QUYcZ3XJVRXWa09Fd_\CW8JI](R_?
7XVfL@OO&H&PfAY7J6DAW1W6O&CM5V+[[L8=88U[eeY4-ED0:1DMLeS0/J;R4f6Y
Q\GJ<34J8VPVF41BRW&O_NER1P9#8CHb4Ab_9Y+;N9R2b#3Z>Uce9/3\]fWT>2M^
;\A_]BB+GfAS#B41^C0edBF?/-d@TQ&3_#]/<.Q@R)>EM1Zd[X].M@D[X6;,Hc1[
X5>:Ta:+HSF?X^c4eDIZC>M:9M#UF&?Q9\?YK7?U2?ZEG$
`endprotected
